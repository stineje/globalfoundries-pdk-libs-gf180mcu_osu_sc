VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffn_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffn_1 ;
  SIZE 14.250 BY 8.300 ;
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.900 3.900 2.400 3.950 ;
        RECT 1.750 3.600 2.550 3.900 ;
        RECT 1.900 3.550 2.400 3.600 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.550 3.250 9.950 3.300 ;
        RECT 9.500 2.950 10.000 3.250 ;
        RECT 9.550 2.900 9.950 2.950 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.450 5.200 13.850 5.250 ;
        RECT 13.400 4.900 13.900 5.200 ;
        RECT 13.450 4.850 13.850 4.900 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 0.765000 ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.700 4.550 13.100 4.600 ;
        RECT 12.650 4.250 13.150 4.550 ;
        RECT 12.700 4.200 13.100 4.250 ;
    END
  END QN
  PIN VDD
    ANTENNADIFFAREA 8.642501 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 14.250 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 14.250 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 4.450 5.550 4.700 7.600 ;
        RECT 7.250 6.300 7.500 7.600 ;
        RECT 9.950 5.550 10.350 7.600 ;
        RECT 12.550 5.550 12.800 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 6.102500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 4.450 0.700 4.700 1.500 ;
        RECT 7.250 0.700 7.500 1.900 ;
        RECT 9.950 0.700 10.350 1.550 ;
        RECT 12.550 0.700 12.800 1.900 ;
        RECT 0.000 0.000 14.250 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.700 0.800 7.250 ;
        RECT 3.050 5.300 3.300 7.250 ;
        RECT 5.850 6.300 6.100 7.250 ;
        RECT 1.400 5.050 3.300 5.300 ;
        RECT 4.950 6.050 6.100 6.300 ;
        RECT 8.100 6.050 8.350 7.250 ;
        RECT 1.400 4.550 1.650 5.050 ;
        RECT 4.050 4.900 4.550 5.200 ;
        RECT 1.050 4.250 1.650 4.550 ;
        RECT 2.600 4.250 3.100 4.550 ;
        RECT 0.500 2.200 0.800 2.700 ;
        RECT 1.400 2.600 1.650 4.250 ;
        RECT 2.700 4.200 3.000 4.250 ;
        RECT 1.900 3.600 2.400 3.900 ;
        RECT 4.150 2.600 4.450 4.900 ;
        RECT 4.950 3.800 5.200 6.050 ;
        RECT 8.100 5.750 8.400 6.050 ;
        RECT 9.100 5.800 9.350 7.250 ;
        RECT 6.000 5.550 8.400 5.750 ;
        RECT 8.950 5.550 9.350 5.800 ;
        RECT 6.000 5.450 8.350 5.550 ;
        RECT 6.000 5.200 6.300 5.450 ;
        RECT 5.900 4.900 6.400 5.200 ;
        RECT 6.700 4.900 7.200 5.200 ;
        RECT 8.100 5.100 8.350 5.450 ;
        RECT 4.900 3.550 5.200 3.800 ;
        RECT 5.500 4.250 6.550 4.550 ;
        RECT 1.400 2.350 2.400 2.600 ;
        RECT 0.550 1.050 0.800 2.200 ;
        RECT 2.000 1.900 2.400 2.350 ;
        RECT 4.050 2.300 4.550 2.600 ;
        RECT 4.900 1.950 5.150 3.550 ;
        RECT 5.500 2.550 5.800 4.250 ;
        RECT 6.800 3.900 7.100 4.900 ;
        RECT 8.100 4.850 8.700 5.100 ;
        RECT 7.650 4.250 8.150 4.550 ;
        RECT 8.400 3.900 8.700 4.850 ;
        RECT 6.750 3.600 7.250 3.900 ;
        RECT 8.100 3.650 8.700 3.900 ;
        RECT 5.400 2.250 5.900 2.550 ;
        RECT 2.000 1.650 3.300 1.900 ;
        RECT 4.900 1.700 6.250 1.950 ;
        RECT 3.050 1.050 3.300 1.650 ;
        RECT 5.850 1.650 6.250 1.700 ;
        RECT 5.850 1.050 6.100 1.650 ;
        RECT 8.100 1.050 8.350 3.650 ;
        RECT 8.950 1.950 9.250 5.550 ;
        RECT 10.300 5.200 10.600 5.300 ;
        RECT 10.200 4.900 10.700 5.200 ;
        RECT 9.600 3.250 9.900 3.350 ;
        RECT 9.500 2.950 10.000 3.250 ;
        RECT 9.600 2.850 9.900 2.950 ;
        RECT 10.300 2.100 10.600 4.900 ;
        RECT 10.950 3.250 11.200 7.250 ;
        RECT 11.700 4.550 11.950 7.250 ;
        RECT 13.400 5.250 13.650 7.250 ;
        RECT 13.400 4.900 13.900 5.250 ;
        RECT 13.400 4.850 13.850 4.900 ;
        RECT 11.700 4.250 13.150 4.550 ;
        RECT 10.950 2.950 12.400 3.250 ;
        RECT 8.950 1.700 9.350 1.950 ;
        RECT 10.200 1.800 10.700 2.100 ;
        RECT 9.100 1.050 9.350 1.700 ;
        RECT 10.950 1.050 11.200 2.950 ;
        RECT 12.800 2.400 13.050 4.250 ;
        RECT 11.700 2.150 13.050 2.400 ;
        RECT 11.700 1.050 11.950 2.150 ;
        RECT 13.400 1.050 13.650 4.850 ;
      LAYER Via1 ;
        RECT 2.700 4.250 3.000 4.550 ;
        RECT 0.500 2.300 0.800 2.600 ;
        RECT 2.000 3.600 2.300 3.900 ;
        RECT 6.800 4.900 7.100 5.200 ;
        RECT 6.150 4.250 6.450 4.550 ;
        RECT 4.150 2.300 4.450 2.600 ;
        RECT 7.750 4.250 8.050 4.550 ;
        RECT 6.850 3.600 7.150 3.900 ;
        RECT 8.950 4.250 9.250 4.550 ;
        RECT 9.600 2.950 9.900 3.250 ;
        RECT 13.500 4.900 13.800 5.200 ;
        RECT 12.750 4.250 13.050 4.550 ;
        RECT 12.000 2.950 12.300 3.250 ;
        RECT 10.300 1.800 10.600 2.100 ;
      LAYER Metal2 ;
        RECT 6.750 5.200 7.150 5.250 ;
        RECT 6.700 4.900 11.150 5.200 ;
        RECT 6.750 4.850 7.150 4.900 ;
        RECT 2.600 4.550 3.050 4.600 ;
        RECT 6.050 4.550 6.550 4.600 ;
        RECT 7.700 4.550 8.100 4.600 ;
        RECT 8.900 4.550 9.300 4.600 ;
        RECT 2.600 4.250 9.350 4.550 ;
        RECT 2.600 4.200 3.050 4.250 ;
        RECT 6.050 4.200 6.550 4.250 ;
        RECT 7.700 4.200 8.100 4.250 ;
        RECT 8.900 4.200 9.300 4.250 ;
        RECT 6.800 3.900 7.200 3.950 ;
        RECT 6.750 3.600 7.250 3.900 ;
        RECT 6.800 3.550 7.200 3.600 ;
        RECT 10.850 3.250 11.150 4.900 ;
        RECT 11.950 3.250 12.350 3.300 ;
        RECT 10.850 2.950 12.400 3.250 ;
        RECT 11.950 2.900 12.350 2.950 ;
        RECT 0.450 2.600 0.850 2.650 ;
        RECT 4.100 2.600 4.500 2.650 ;
        RECT 0.400 2.300 4.550 2.600 ;
        RECT 0.450 2.250 0.850 2.300 ;
        RECT 4.100 2.250 4.500 2.300 ;
        RECT 10.250 2.100 10.650 2.150 ;
        RECT 5.800 1.950 6.200 2.000 ;
        RECT 9.500 1.950 10.700 2.100 ;
        RECT 5.750 1.800 10.700 1.950 ;
        RECT 5.750 1.750 10.650 1.800 ;
        RECT 5.750 1.650 9.900 1.750 ;
        RECT 5.800 1.600 6.200 1.650 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffn_1


MACRO gf180mcu_osu_sc_gp12t3v3__addh_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addh_1 ;
  SIZE 8.100 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.500 3.900 2.000 3.950 ;
        RECT 3.900 3.900 4.400 3.950 ;
        RECT 1.500 3.600 4.400 3.900 ;
        RECT 1.500 3.550 2.000 3.600 ;
        RECT 3.900 3.550 4.400 3.600 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.350 3.250 2.850 3.300 ;
        RECT 5.200 3.250 5.700 3.300 ;
        RECT 2.350 2.950 5.700 3.250 ;
        RECT 2.350 2.900 2.850 2.950 ;
        RECT 5.200 2.900 5.700 2.950 ;
    END
  END B
  PIN SUM
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.200 4.850 7.700 5.250 ;
    END
  END SUM
  PIN CO
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 2.250 0.900 2.650 ;
    END
  END CO
  PIN VDD
    ANTENNADIFFAREA 5.595000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 8.100 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 8.100 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
        RECT 3.850 5.550 4.100 7.600 ;
        RECT 6.400 5.550 6.650 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.960000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 6.400 0.700 6.650 1.900 ;
        RECT 0.000 0.000 8.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.600 0.800 7.250 ;
        RECT 2.250 5.200 2.500 7.250 ;
        RECT 1.050 4.900 3.500 5.200 ;
        RECT 1.500 3.600 2.000 3.900 ;
        RECT 2.350 2.950 2.850 3.250 ;
        RECT 0.400 2.300 0.900 2.600 ;
        RECT 0.550 1.050 0.800 2.300 ;
        RECT 3.100 1.050 3.350 4.900 ;
        RECT 5.550 3.900 5.800 7.250 ;
        RECT 7.250 5.250 7.500 7.250 ;
        RECT 7.250 5.200 7.600 5.250 ;
        RECT 6.050 4.900 6.550 5.200 ;
        RECT 7.200 4.900 7.700 5.200 ;
        RECT 7.250 4.850 7.600 4.900 ;
        RECT 3.900 3.600 4.400 3.900 ;
        RECT 5.550 3.850 7.000 3.900 ;
        RECT 4.700 3.600 7.000 3.850 ;
        RECT 3.850 1.200 4.100 2.000 ;
        RECT 4.700 1.450 4.950 3.600 ;
        RECT 5.200 2.950 5.700 3.250 ;
        RECT 5.550 1.200 5.800 2.000 ;
        RECT 3.850 0.950 5.800 1.200 ;
        RECT 7.250 1.050 7.500 4.850 ;
      LAYER Via1 ;
        RECT 3.100 4.900 3.400 5.200 ;
        RECT 1.600 3.600 1.900 3.900 ;
        RECT 2.450 2.950 2.750 3.250 ;
        RECT 0.500 2.300 0.800 2.600 ;
        RECT 6.150 4.900 6.450 5.200 ;
        RECT 7.300 4.900 7.600 5.200 ;
        RECT 4.000 3.600 4.300 3.900 ;
        RECT 5.300 2.950 5.600 3.250 ;
      LAYER Metal2 ;
        RECT 3.000 5.200 3.500 5.250 ;
        RECT 6.050 5.200 6.550 5.250 ;
        RECT 3.000 4.900 6.550 5.200 ;
        RECT 3.000 4.850 3.500 4.900 ;
        RECT 6.050 4.850 6.550 4.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addh_1


MACRO gf180mcu_osu_sc_gp12t3v3__tieh
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tieh ;
  SIZE 2.200 BY 8.300 ;
  PIN Y
    ANTENNADIFFAREA 0.850000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 4.850 1.800 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 2.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 2.200 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.762500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 5.200 1.650 7.250 ;
        RECT 1.300 4.900 1.800 5.200 ;
        RECT 1.400 4.850 1.650 4.900 ;
        RECT 1.150 2.300 1.650 2.550 ;
        RECT 1.400 1.050 1.650 2.300 ;
      LAYER Via1 ;
        RECT 1.400 4.900 1.700 5.200 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tieh


MACRO gf180mcu_osu_sc_gp12t3v3__fill_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_8 ;
  SIZE 0.900 BY 8.300 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.600 0.800 8.300 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 0.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 5.100 0.800 8.300 ;
  END
END gf180mcu_osu_sc_gp12t3v3__fill_8


MACRO gf180mcu_osu_sc_gp12t3v3__xnor2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__xnor2_1 ;
  SIZE 6.200 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.650 3.950 3.950 4.000 ;
        RECT 3.600 3.550 4.000 3.950 ;
        RECT 1.350 2.650 1.650 2.700 ;
        RECT 1.300 2.250 1.700 2.650 ;
        RECT 1.350 1.300 1.650 2.250 ;
        RECT 3.650 1.300 3.950 3.550 ;
        RECT 1.350 1.000 3.950 1.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 4.450 2.650 4.750 2.700 ;
        RECT 4.400 2.600 4.800 2.650 ;
        RECT 4.350 2.300 4.850 2.600 ;
        RECT 4.400 2.250 4.800 2.300 ;
        RECT 4.450 2.200 4.750 2.250 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 2.192500 ;
    PORT
      LAYER Metal2 ;
        RECT 2.900 5.900 3.200 6.050 ;
        RECT 2.850 5.500 3.250 5.900 ;
        RECT 2.900 2.000 3.200 5.500 ;
        RECT 2.800 1.600 3.300 2.000 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.557500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 6.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 6.200 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 4.500 5.550 4.750 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.622500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 4.500 0.700 4.750 1.900 ;
        RECT 0.000 0.000 6.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.900 0.800 7.250 ;
        RECT 2.950 5.950 3.200 7.250 ;
        RECT 2.900 5.400 3.200 5.950 ;
        RECT 5.350 4.550 5.600 7.250 ;
        RECT 2.550 4.250 5.600 4.550 ;
        RECT 0.550 3.600 3.300 3.900 ;
        RECT 3.550 3.600 4.050 3.900 ;
        RECT 0.550 1.050 0.800 3.600 ;
        RECT 3.000 2.600 3.300 3.600 ;
        RECT 1.250 2.300 1.750 2.600 ;
        RECT 2.900 2.300 3.400 2.600 ;
        RECT 4.350 2.300 4.850 2.600 ;
        RECT 2.900 1.500 3.200 2.050 ;
        RECT 2.950 1.050 3.200 1.500 ;
        RECT 5.350 1.050 5.600 4.250 ;
      LAYER Via1 ;
        RECT 2.900 5.550 3.200 5.850 ;
        RECT 3.650 3.600 3.950 3.900 ;
        RECT 1.350 2.300 1.650 2.600 ;
        RECT 4.450 2.300 4.750 2.600 ;
        RECT 2.900 1.650 3.200 1.950 ;
  END
END gf180mcu_osu_sc_gp12t3v3__xnor2_1


MACRO gf180mcu_osu_sc_gp12t3v3__aoi22_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi22_1 ;
  SIZE 5.350 BY 8.300 ;
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.600 4.200 2.100 4.600 ;
    END
  END A1
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 3.550 1.100 3.950 ;
    END
  END A0
  PIN B0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.350 3.550 2.850 3.950 ;
    END
  END B0
  PIN B1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.300 4.200 3.800 4.600 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 3.000 6.500 3.500 6.550 ;
        RECT 4.350 6.500 4.850 6.550 ;
        RECT 3.000 6.200 4.850 6.500 ;
        RECT 3.000 6.150 3.500 6.200 ;
        RECT 4.350 6.150 4.850 6.200 ;
        RECT 4.300 4.850 4.800 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.285000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 5.350 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 5.350 8.300 ;
        RECT 1.400 6.300 1.650 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.200000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 0.700 0.950 1.900 ;
        RECT 3.500 0.700 3.750 1.900 ;
        RECT 0.000 0.000 5.350 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 5.950 0.800 7.250 ;
        RECT 2.250 5.950 2.500 7.250 ;
        RECT 3.100 6.500 3.350 7.250 ;
        RECT 3.000 6.200 3.500 6.500 ;
        RECT 3.950 5.950 4.200 7.250 ;
        RECT 0.550 5.700 4.200 5.950 ;
        RECT 4.450 6.100 4.750 6.600 ;
        RECT 4.450 5.200 4.700 6.100 ;
        RECT 4.300 4.900 4.800 5.200 ;
        RECT 1.600 4.250 2.100 4.550 ;
        RECT 3.300 4.250 3.800 4.550 ;
        RECT 0.600 3.600 1.100 3.900 ;
        RECT 2.350 3.600 2.850 3.900 ;
        RECT 4.400 3.350 4.650 4.900 ;
        RECT 2.100 3.100 4.650 3.350 ;
        RECT 2.100 1.050 2.350 3.100 ;
      LAYER Via1 ;
        RECT 3.100 6.200 3.400 6.500 ;
        RECT 4.450 6.200 4.750 6.500 ;
        RECT 4.400 4.900 4.700 5.200 ;
        RECT 1.700 4.250 2.000 4.550 ;
        RECT 3.400 4.250 3.700 4.550 ;
        RECT 0.700 3.600 1.000 3.900 ;
        RECT 2.450 3.600 2.750 3.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi22_1


MACRO gf180mcu_osu_sc_gp12t3v3__dffsr_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsr_1 ;
  SIZE 18.700 BY 8.300 ;
  PIN D
    ANTENNAGATEAREA 0.690000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.950 3.550 6.450 3.950 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.295000 ;
    PORT
      LAYER Metal2 ;
        RECT 6.650 4.550 7.100 4.600 ;
        RECT 10.100 4.550 10.600 4.600 ;
        RECT 11.750 4.550 12.150 4.600 ;
        RECT 6.650 4.250 12.200 4.550 ;
        RECT 6.650 4.200 7.100 4.250 ;
        RECT 10.100 4.200 10.600 4.250 ;
        RECT 11.750 4.200 12.150 4.250 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.950 5.200 18.350 5.250 ;
        RECT 17.900 4.900 18.400 5.200 ;
        RECT 17.950 4.850 18.350 4.900 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 0.765000 ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.200 4.550 17.600 4.600 ;
        RECT 17.150 4.250 17.650 4.550 ;
        RECT 17.200 4.200 17.600 4.250 ;
    END
  END QN
  PIN R
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.550 4.850 1.050 5.250 ;
    END
  END R
  PIN VDD
    ANTENNADIFFAREA 11.437501 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 18.700 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 18.700 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 3.850 6.300 4.100 7.600 ;
        RECT 5.450 5.550 5.700 7.600 ;
        RECT 8.500 5.550 8.750 7.600 ;
        RECT 11.300 6.300 11.550 7.600 ;
        RECT 13.750 6.800 14.000 7.600 ;
        RECT 17.050 5.550 17.300 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.940001 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.300 0.700 2.550 1.900 ;
        RECT 4.550 0.700 4.800 1.900 ;
        RECT 5.450 0.700 5.700 1.900 ;
        RECT 8.500 0.700 8.750 1.500 ;
        RECT 11.300 0.700 11.550 1.900 ;
        RECT 13.050 0.700 13.300 1.900 ;
        RECT 15.300 0.700 15.550 1.900 ;
        RECT 17.050 0.700 17.300 1.900 ;
        RECT 0.000 0.000 18.700 0.700 ;
    END
  END VSS
  PIN S
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.500 5.550 14.350 5.850 ;
        RECT 3.500 4.600 3.800 5.550 ;
        RECT 14.050 4.600 14.350 5.550 ;
        RECT 3.400 4.200 3.900 4.600 ;
        RECT 13.950 4.200 14.450 4.600 ;
    END
  END S
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.900 1.050 5.200 ;
        RECT 1.400 2.600 1.650 7.250 ;
        RECT 2.150 2.850 2.400 7.250 ;
        RECT 3.000 6.050 3.250 7.250 ;
        RECT 4.700 6.050 4.950 7.250 ;
        RECT 3.000 5.800 4.950 6.050 ;
        RECT 7.100 5.300 7.350 7.250 ;
        RECT 9.900 6.300 10.150 7.250 ;
        RECT 5.450 5.050 7.350 5.300 ;
        RECT 9.000 6.050 10.150 6.300 ;
        RECT 3.400 4.250 3.900 4.550 ;
        RECT 5.450 3.900 5.700 5.050 ;
        RECT 8.100 4.900 8.600 5.200 ;
        RECT 6.650 4.250 7.650 4.550 ;
        RECT 6.750 4.200 7.050 4.250 ;
        RECT 2.650 3.600 3.150 3.900 ;
        RECT 4.400 3.600 5.700 3.900 ;
        RECT 5.950 3.600 6.450 3.900 ;
        RECT 2.150 2.600 3.400 2.850 ;
        RECT 4.500 2.600 4.750 2.650 ;
        RECT 5.450 2.600 5.700 3.600 ;
        RECT 1.300 2.300 1.800 2.600 ;
        RECT 3.150 2.300 4.900 2.600 ;
        RECT 5.450 2.350 6.450 2.600 ;
        RECT 7.350 2.450 7.650 4.250 ;
        RECT 8.200 2.600 8.500 4.900 ;
        RECT 9.000 3.800 9.250 6.050 ;
        RECT 10.100 5.250 10.400 5.350 ;
        RECT 10.000 4.950 10.500 5.250 ;
        RECT 10.100 4.550 10.400 4.950 ;
        RECT 10.750 4.900 11.250 5.200 ;
        RECT 12.150 5.100 12.400 7.250 ;
        RECT 12.900 6.550 13.150 7.250 ;
        RECT 14.600 6.550 14.850 7.250 ;
        RECT 12.900 6.300 14.850 6.550 ;
        RECT 13.050 5.200 13.350 5.300 ;
        RECT 15.450 5.200 15.700 7.250 ;
        RECT 8.950 3.550 9.250 3.800 ;
        RECT 9.550 4.250 10.600 4.550 ;
        RECT 1.400 2.250 1.700 2.300 ;
        RECT 1.400 1.050 1.650 2.250 ;
        RECT 3.150 1.050 3.400 2.300 ;
        RECT 4.500 2.250 4.750 2.300 ;
        RECT 6.050 1.900 6.450 2.350 ;
        RECT 7.250 2.150 7.750 2.450 ;
        RECT 8.100 2.300 8.600 2.600 ;
        RECT 8.950 1.950 9.200 3.550 ;
        RECT 9.550 2.550 9.850 4.250 ;
        RECT 10.850 3.900 11.150 4.900 ;
        RECT 12.150 4.850 12.700 5.100 ;
        RECT 11.700 4.250 12.200 4.550 ;
        RECT 12.450 3.900 12.700 4.850 ;
        RECT 13.050 4.900 15.850 5.200 ;
        RECT 13.050 4.800 13.350 4.900 ;
        RECT 13.950 4.250 14.450 4.550 ;
        RECT 10.800 3.600 11.300 3.900 ;
        RECT 12.150 3.650 12.700 3.900 ;
        RECT 10.100 2.950 10.600 3.250 ;
        RECT 12.150 2.850 12.450 3.650 ;
        RECT 15.450 3.250 15.700 4.900 ;
        RECT 16.200 4.550 16.450 7.250 ;
        RECT 17.900 5.250 18.150 7.250 ;
        RECT 17.900 4.900 18.400 5.250 ;
        RECT 17.900 4.850 18.350 4.900 ;
        RECT 16.200 4.250 17.650 4.550 ;
        RECT 14.450 2.950 16.900 3.250 ;
        RECT 9.450 2.250 9.950 2.550 ;
        RECT 6.050 1.650 7.350 1.900 ;
        RECT 8.950 1.700 10.300 1.950 ;
        RECT 7.100 1.050 7.350 1.650 ;
        RECT 9.900 1.650 10.300 1.700 ;
        RECT 9.900 1.050 10.150 1.650 ;
        RECT 12.150 1.050 12.400 2.850 ;
        RECT 12.950 2.250 13.450 2.550 ;
        RECT 14.450 1.050 14.700 2.950 ;
        RECT 14.950 2.250 15.450 2.550 ;
        RECT 17.300 2.400 17.550 4.250 ;
        RECT 16.200 2.150 17.550 2.400 ;
        RECT 16.200 1.050 16.450 2.150 ;
        RECT 17.900 1.050 18.150 4.850 ;
      LAYER Via1 ;
        RECT 0.650 4.900 0.950 5.200 ;
        RECT 3.500 4.250 3.800 4.550 ;
        RECT 6.750 4.250 7.050 4.550 ;
        RECT 2.750 3.600 3.050 3.900 ;
        RECT 4.500 3.600 4.800 3.900 ;
        RECT 6.050 3.600 6.350 3.900 ;
        RECT 1.400 2.300 1.700 2.600 ;
        RECT 4.500 2.300 4.800 2.600 ;
        RECT 10.850 4.900 11.150 5.200 ;
        RECT 10.200 4.250 10.500 4.550 ;
        RECT 8.200 2.300 8.500 2.600 ;
        RECT 11.800 4.250 12.100 4.550 ;
        RECT 15.450 4.900 15.750 5.200 ;
        RECT 14.050 4.250 14.350 4.550 ;
        RECT 10.900 3.600 11.200 3.900 ;
        RECT 18.000 4.900 18.300 5.200 ;
        RECT 17.250 4.250 17.550 4.550 ;
        RECT 10.200 2.950 10.500 3.250 ;
        RECT 12.150 2.950 12.450 3.250 ;
        RECT 16.500 2.950 16.800 3.250 ;
        RECT 13.050 2.250 13.350 2.550 ;
        RECT 15.050 2.250 15.350 2.550 ;
      LAYER Metal2 ;
        RECT 10.800 5.200 11.200 5.250 ;
        RECT 13.000 5.200 13.400 5.250 ;
        RECT 10.750 4.900 13.450 5.200 ;
        RECT 10.800 4.850 11.200 4.900 ;
        RECT 13.000 4.850 13.400 4.900 ;
        RECT 15.350 4.850 15.850 5.250 ;
        RECT 2.650 3.550 3.150 3.950 ;
        RECT 4.400 3.550 4.900 3.950 ;
        RECT 10.850 3.900 11.250 3.950 ;
        RECT 10.800 3.600 11.300 3.900 ;
        RECT 10.850 3.550 11.250 3.600 ;
        RECT 1.300 2.600 1.800 2.650 ;
        RECT 2.750 2.600 3.050 3.550 ;
        RECT 10.150 3.250 10.550 3.300 ;
        RECT 12.100 3.250 12.500 3.300 ;
        RECT 16.450 3.250 16.850 3.300 ;
        RECT 10.100 2.950 12.600 3.250 ;
        RECT 16.100 2.950 16.900 3.250 ;
        RECT 10.150 2.900 10.550 2.950 ;
        RECT 12.100 2.900 12.500 2.950 ;
        RECT 16.450 2.900 16.850 2.950 ;
        RECT 1.300 2.300 3.050 2.600 ;
        RECT 1.300 2.250 1.800 2.300 ;
        RECT 2.750 1.300 3.050 2.300 ;
        RECT 4.400 2.600 4.900 2.650 ;
        RECT 8.150 2.600 8.550 2.650 ;
        RECT 4.400 2.300 8.600 2.600 ;
        RECT 4.400 2.250 4.900 2.300 ;
        RECT 8.150 2.250 8.550 2.300 ;
        RECT 12.950 2.200 13.450 2.600 ;
        RECT 14.850 2.200 15.450 2.600 ;
        RECT 9.850 1.950 10.250 2.000 ;
        RECT 12.950 1.950 13.350 2.200 ;
        RECT 9.800 1.650 13.350 1.950 ;
        RECT 9.850 1.600 10.250 1.650 ;
        RECT 14.850 1.300 15.150 2.200 ;
        RECT 2.750 1.000 15.150 1.300 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsr_1


MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_8 ;
  SIZE 8.150 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 6.120000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 3.550 0.900 3.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 5.610001 ;
    PORT
      LAYER Metal2 ;
        RECT 6.350 4.450 6.850 4.850 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 6.530001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 8.150 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 8.150 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
        RECT 3.950 5.550 4.200 7.600 ;
        RECT 5.650 5.550 5.900 7.600 ;
        RECT 7.350 5.550 7.600 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.277500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 5.650 0.700 5.900 1.900 ;
        RECT 7.350 0.700 7.600 1.900 ;
        RECT 0.000 0.000 8.150 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.800 1.650 7.250 ;
        RECT 3.100 4.800 3.350 7.250 ;
        RECT 4.800 4.800 5.050 7.250 ;
        RECT 6.500 4.800 6.750 7.250 ;
        RECT 1.400 4.550 6.750 4.800 ;
        RECT 0.400 3.600 0.900 3.900 ;
        RECT 1.400 2.400 1.650 4.550 ;
        RECT 3.100 2.400 3.350 4.550 ;
        RECT 4.800 2.400 5.050 4.550 ;
        RECT 6.350 4.450 6.750 4.550 ;
        RECT 6.500 2.400 6.750 4.450 ;
        RECT 1.400 2.150 6.750 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
        RECT 4.800 1.050 5.050 2.150 ;
        RECT 6.500 1.050 6.750 2.150 ;
      LAYER Via1 ;
        RECT 0.500 3.600 0.800 3.900 ;
        RECT 6.450 4.500 6.750 4.800 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkinv_8


MACRO gf180mcu_osu_sc_gp12t3v3__inv_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_16 ;
  SIZE 15.000 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 12.240001 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 3.550 0.900 3.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 11.220001 ;
    PORT
      LAYER Metal2 ;
        RECT 13.150 4.200 13.650 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 12.295001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 15.000 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 15.000 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
        RECT 3.950 5.550 4.200 7.600 ;
        RECT 5.650 5.550 5.900 7.600 ;
        RECT 7.350 5.550 7.600 7.600 ;
        RECT 9.050 5.550 9.300 7.600 ;
        RECT 10.750 5.550 11.000 7.600 ;
        RECT 12.450 5.550 12.700 7.600 ;
        RECT 14.150 5.550 14.400 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.172501 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 5.650 0.700 5.900 1.900 ;
        RECT 7.350 0.700 7.600 1.900 ;
        RECT 9.050 0.700 9.300 1.900 ;
        RECT 10.750 0.700 11.000 1.900 ;
        RECT 12.450 0.700 12.700 1.900 ;
        RECT 14.150 0.700 14.400 1.900 ;
        RECT 0.000 0.000 15.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.800 1.650 7.250 ;
        RECT 3.100 4.800 3.350 7.250 ;
        RECT 4.800 4.800 5.050 7.250 ;
        RECT 6.500 4.800 6.750 7.250 ;
        RECT 8.200 4.800 8.450 7.250 ;
        RECT 9.900 4.800 10.150 7.250 ;
        RECT 11.600 4.800 11.850 7.250 ;
        RECT 13.300 4.800 13.550 7.250 ;
        RECT 1.400 4.550 13.550 4.800 ;
        RECT 0.400 3.600 0.900 3.900 ;
        RECT 1.400 2.400 1.650 4.550 ;
        RECT 3.100 2.400 3.350 4.550 ;
        RECT 4.800 2.400 5.050 4.550 ;
        RECT 6.500 2.400 6.750 4.550 ;
        RECT 8.200 2.400 8.450 4.550 ;
        RECT 9.900 2.400 10.150 4.550 ;
        RECT 11.600 2.400 11.850 4.550 ;
        RECT 13.150 4.200 13.550 4.550 ;
        RECT 13.300 2.400 13.550 4.200 ;
        RECT 1.400 2.150 13.550 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
        RECT 4.800 1.050 5.050 2.150 ;
        RECT 6.500 1.050 6.750 2.150 ;
        RECT 8.200 1.050 8.450 2.150 ;
        RECT 9.900 1.050 10.150 2.150 ;
        RECT 11.600 1.050 11.850 2.150 ;
        RECT 13.300 1.050 13.550 2.150 ;
      LAYER Via1 ;
        RECT 0.500 3.600 0.800 3.900 ;
        RECT 13.250 4.250 13.550 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__inv_16


MACRO gf180mcu_osu_sc_gp12t3v3__oai22_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai22_1 ;
  SIZE 5.300 BY 8.300 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.450 3.550 0.950 3.950 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.450 4.200 1.950 4.600 ;
    END
  END A1
  PIN B0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.200 3.550 2.700 3.950 ;
    END
  END B0
  PIN B1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 3.550 3.650 3.950 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 4.300 4.200 4.800 4.600 ;
        RECT 2.950 1.300 3.450 1.350 ;
        RECT 4.350 1.300 4.750 1.450 ;
        RECT 2.950 1.000 4.750 1.300 ;
        RECT 2.950 0.950 3.450 1.000 ;
        RECT 4.350 0.950 4.750 1.000 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.050000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 5.300 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 5.300 8.300 ;
        RECT 0.650 5.550 0.900 7.600 ;
        RECT 3.500 5.550 3.750 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.817500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 0.700 1.600 1.700 ;
        RECT 0.000 0.000 5.300 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.100 5.300 2.350 7.250 ;
        RECT 2.100 5.000 4.650 5.300 ;
        RECT 4.400 4.550 4.650 5.000 ;
        RECT 1.450 4.250 1.950 4.550 ;
        RECT 4.300 4.250 4.800 4.550 ;
        RECT 0.450 3.600 0.950 3.900 ;
        RECT 2.200 3.600 2.700 3.900 ;
        RECT 3.150 3.600 3.650 3.900 ;
        RECT 0.500 1.950 4.150 2.200 ;
        RECT 0.500 1.050 0.750 1.950 ;
        RECT 2.200 1.050 2.450 1.950 ;
        RECT 3.050 1.300 3.300 1.700 ;
        RECT 2.950 1.000 3.450 1.300 ;
        RECT 3.900 1.050 4.150 1.950 ;
        RECT 4.400 1.450 4.650 4.250 ;
        RECT 4.400 0.950 4.700 1.450 ;
      LAYER Via1 ;
        RECT 1.550 4.250 1.850 4.550 ;
        RECT 4.400 4.250 4.700 4.550 ;
        RECT 0.550 3.600 0.850 3.900 ;
        RECT 2.300 3.600 2.600 3.900 ;
        RECT 3.250 3.600 3.550 3.900 ;
        RECT 3.050 1.000 3.350 1.300 ;
        RECT 4.400 1.050 4.700 1.350 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai22_1


MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_1 ;
  SIZE 2.200 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.550 4.850 1.050 5.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 3.550 1.800 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 2.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 2.200 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.762500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.900 1.050 5.200 ;
        RECT 1.400 3.900 1.650 7.250 ;
        RECT 1.300 3.600 1.800 3.900 ;
        RECT 1.400 1.050 1.650 3.600 ;
      LAYER Via1 ;
        RECT 0.650 4.900 0.950 5.200 ;
        RECT 1.400 3.600 1.700 3.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkinv_1


MACRO gf180mcu_osu_sc_gp12t3v3__addf_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addf_1 ;
  SIZE 14.000 BY 8.350 ;
  PIN A
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.650 3.900 1.050 3.950 ;
        RECT 4.650 3.900 5.050 3.950 ;
        RECT 8.750 3.900 9.150 3.950 ;
        RECT 0.600 3.600 9.200 3.900 ;
        RECT 0.650 3.550 1.050 3.600 ;
        RECT 4.650 3.550 5.050 3.600 ;
        RECT 8.750 3.550 9.150 3.600 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.550 4.550 1.950 4.600 ;
        RECT 3.650 4.550 4.050 4.600 ;
        RECT 5.800 4.550 6.200 4.600 ;
        RECT 9.600 4.550 10.000 4.600 ;
        RECT 1.500 4.250 4.100 4.550 ;
        RECT 5.750 4.250 10.050 4.550 ;
        RECT 1.550 4.200 1.950 4.250 ;
        RECT 3.650 4.200 4.050 4.250 ;
        RECT 5.800 4.200 6.200 4.250 ;
        RECT 9.600 4.200 10.000 4.250 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA 2.295000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.400 3.250 2.800 3.300 ;
        RECT 2.350 2.950 2.850 3.250 ;
        RECT 2.400 2.900 2.800 2.950 ;
        RECT 2.450 2.600 2.750 2.900 ;
        RECT 6.700 2.600 7.100 2.650 ;
        RECT 10.100 2.600 10.500 2.650 ;
        RECT 2.450 2.300 10.550 2.600 ;
        RECT 6.700 2.250 7.100 2.300 ;
        RECT 10.100 2.250 10.500 2.300 ;
        RECT 6.750 2.200 7.050 2.250 ;
        RECT 10.150 2.200 10.450 2.250 ;
    END
  END CI
  PIN SUM
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.550 4.550 11.950 4.600 ;
        RECT 11.500 4.250 12.000 4.550 ;
        RECT 11.550 4.200 11.950 4.250 ;
    END
  END SUM
  PIN CO
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.300 3.250 13.700 3.300 ;
        RECT 13.250 2.950 13.750 3.250 ;
        RECT 13.300 2.900 13.700 2.950 ;
    END
  END CO
  PIN VSS
    ANTENNADIFFAREA 6.007501 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.550 ;
        RECT 10.750 0.700 11.000 1.900 ;
        RECT 12.350 0.700 12.600 1.900 ;
        RECT 0.000 0.000 14.000 0.700 ;
    END
  END VSS
  PIN VDD
    ANTENNADIFFAREA 8.302501 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 14.000 8.350 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 14.000 8.350 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 4.800 5.550 5.050 7.600 ;
        RECT 6.500 5.550 6.750 7.600 ;
        RECT 10.750 5.550 11.000 7.600 ;
        RECT 12.350 5.550 12.600 7.600 ;
    END
  END VDD
  OBS
      LAYER Metal1 ;
        RECT 0.550 5.300 0.800 7.250 ;
        RECT 2.250 5.300 2.500 7.250 ;
        RECT 0.550 5.050 2.500 5.300 ;
        RECT 1.500 4.250 2.000 4.550 ;
        RECT 0.600 3.600 1.100 3.900 ;
        RECT 3.100 3.250 3.350 7.250 ;
        RECT 5.650 5.300 5.900 7.250 ;
        RECT 7.350 5.300 7.600 7.250 ;
        RECT 5.650 5.050 7.600 5.300 ;
        RECT 3.600 4.250 6.250 4.550 ;
        RECT 4.600 3.600 5.100 3.900 ;
        RECT 8.200 3.250 8.450 7.250 ;
        RECT 11.600 4.550 11.850 7.250 ;
        RECT 9.550 4.250 10.050 4.550 ;
        RECT 11.600 4.250 12.000 4.550 ;
        RECT 8.700 3.600 9.200 3.900 ;
        RECT 2.350 2.950 2.850 3.250 ;
        RECT 3.100 2.950 7.950 3.250 ;
        RECT 8.200 2.950 11.350 3.250 ;
        RECT 0.550 2.150 2.500 2.400 ;
        RECT 0.550 1.050 0.800 2.150 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.100 1.050 3.350 2.950 ;
        RECT 6.650 2.300 7.150 2.600 ;
        RECT 5.650 1.800 7.600 2.050 ;
        RECT 5.650 1.050 5.900 1.800 ;
        RECT 7.350 1.050 7.600 1.800 ;
        RECT 8.200 1.050 8.450 2.950 ;
        RECT 10.050 2.300 10.550 2.600 ;
        RECT 11.600 1.050 11.850 4.250 ;
        RECT 13.200 3.300 13.450 7.250 ;
        RECT 13.200 3.250 13.600 3.300 ;
        RECT 12.450 2.950 12.950 3.250 ;
        RECT 13.200 2.950 13.750 3.250 ;
        RECT 13.200 2.900 13.600 2.950 ;
        RECT 13.200 1.050 13.450 2.900 ;
      LAYER Via1 ;
        RECT 1.600 4.250 1.900 4.550 ;
        RECT 0.700 3.600 1.000 3.900 ;
        RECT 3.700 4.250 4.000 4.550 ;
        RECT 5.850 4.250 6.150 4.550 ;
        RECT 4.700 3.600 5.000 3.900 ;
        RECT 9.650 4.250 9.950 4.550 ;
        RECT 8.800 3.600 9.100 3.900 ;
        RECT 2.450 2.950 2.750 3.250 ;
        RECT 7.550 2.950 7.850 3.250 ;
        RECT 6.750 2.300 7.050 2.600 ;
        RECT 10.150 2.300 10.450 2.600 ;
        RECT 12.550 2.950 12.850 3.250 ;
        RECT 13.350 2.950 13.650 3.250 ;
      LAYER Metal2 ;
        RECT 7.500 3.250 7.900 3.300 ;
        RECT 12.500 3.250 12.900 3.300 ;
        RECT 7.450 2.950 12.950 3.250 ;
        RECT 7.500 2.900 7.900 2.950 ;
        RECT 12.500 2.900 12.900 2.950 ;
        RECT 12.550 2.850 12.850 2.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addf_1


MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_8 ;
  SIZE 9.000 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 5.610001 ;
    PORT
      LAYER Metal2 ;
        RECT 7.250 5.250 7.750 5.300 ;
        RECT 7.200 4.950 7.750 5.250 ;
        RECT 7.250 4.900 7.750 4.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 6.615000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 9.000 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 9.000 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
        RECT 4.800 5.550 5.050 7.600 ;
        RECT 6.500 5.550 6.750 7.600 ;
        RECT 8.200 5.550 8.450 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.900 ;
        RECT 8.200 0.700 8.450 1.900 ;
        RECT 0.000 0.000 9.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.250 2.500 7.250 ;
        RECT 3.950 5.250 4.200 7.250 ;
        RECT 5.650 5.250 5.900 7.250 ;
        RECT 7.350 5.250 7.600 7.250 ;
        RECT 2.250 4.950 7.750 5.250 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 2.400 2.500 4.950 ;
        RECT 3.950 2.400 4.200 4.950 ;
        RECT 5.650 2.400 5.900 4.950 ;
        RECT 7.350 2.400 7.600 4.950 ;
        RECT 2.250 2.150 7.600 2.400 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
        RECT 5.650 1.050 5.900 2.150 ;
        RECT 7.350 1.050 7.600 2.150 ;
      LAYER Via1 ;
        RECT 7.350 4.950 7.650 5.250 ;
        RECT 1.150 4.250 1.450 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_8


MACRO gf180mcu_osu_sc_gp12t3v3__lshifdown
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifdown ;
  SIZE 5.200 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 2.250 1.100 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 4.250 4.200 4.750 4.600 ;
    END
  END Y
  PIN VDDH
    ANTENNADIFFAREA 1.272500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 2.300 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 2.300 8.300 ;
        RECT 0.550 5.550 0.850 7.600 ;
    END
  END VDDH
  PIN VDD
    ANTENNADIFFAREA 1.272500 ;
    PORT
      LAYER Nwell ;
        RECT 2.900 5.100 5.200 8.300 ;
      LAYER Metal1 ;
        RECT 2.900 7.600 5.200 8.300 ;
        RECT 3.450 5.550 3.750 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.610000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.850 1.900 ;
        RECT 3.450 0.700 3.750 1.900 ;
        RECT 0.000 0.000 5.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.450 5.200 1.750 7.250 ;
        RECT 1.350 4.900 1.850 5.200 ;
        RECT 3.500 4.900 4.000 5.200 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 1.450 1.050 1.750 4.900 ;
        RECT 4.350 4.550 4.650 7.250 ;
        RECT 4.300 4.250 4.700 4.550 ;
        RECT 4.350 1.050 4.650 4.250 ;
      LAYER Via1 ;
        RECT 1.450 4.900 1.750 5.200 ;
        RECT 3.600 4.900 3.900 5.200 ;
        RECT 0.700 2.300 1.000 2.600 ;
        RECT 4.350 4.250 4.650 4.550 ;
      LAYER Metal2 ;
        RECT 1.350 5.200 1.850 5.250 ;
        RECT 3.500 5.200 4.000 5.250 ;
        RECT 1.350 4.900 4.000 5.200 ;
        RECT 1.350 4.850 1.850 4.900 ;
        RECT 3.500 4.850 4.000 4.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifdown


MACRO gf180mcu_osu_sc_gp12t3v3__buf_4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_4 ;
  SIZE 5.600 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.805000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.800 4.950 4.350 5.250 ;
        RECT 3.850 4.850 4.350 4.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 4.070000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 5.600 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 5.600 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
        RECT 4.800 5.550 5.050 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.710000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 0.000 0.000 5.600 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.250 2.500 7.250 ;
        RECT 3.950 5.250 4.200 7.250 ;
        RECT 2.250 5.200 4.200 5.250 ;
        RECT 2.250 4.950 4.350 5.200 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 2.400 2.500 4.950 ;
        RECT 3.850 4.900 4.350 4.950 ;
        RECT 3.950 2.400 4.200 4.900 ;
        RECT 2.250 2.150 4.200 2.400 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
      LAYER Via1 ;
        RECT 1.150 4.250 1.450 4.550 ;
        RECT 3.950 4.900 4.250 5.200 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_4


MACRO gf180mcu_osu_sc_gp12t3v3__dlat_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dlat_1 ;
  SIZE 9.000 BY 8.300 ;
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.850 4.200 2.350 4.600 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.500 4.550 3.900 4.600 ;
        RECT 5.200 4.550 5.700 4.600 ;
        RECT 3.450 4.250 5.700 4.550 ;
        RECT 3.500 4.200 3.900 4.250 ;
        RECT 5.200 4.200 5.700 4.250 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.200 5.200 8.600 5.250 ;
        RECT 8.150 4.900 8.650 5.200 ;
        RECT 8.200 4.850 8.600 4.900 ;
    END
  END Q
  PIN VDD
    ANTENNADIFFAREA 5.167500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 9.000 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 9.000 8.300 ;
        RECT 1.450 6.350 1.700 7.600 ;
        RECT 4.850 5.550 5.100 7.600 ;
        RECT 7.300 5.550 7.550 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.020000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 0.700 1.850 1.900 ;
        RECT 4.700 0.700 5.100 1.900 ;
        RECT 7.300 0.700 7.550 1.900 ;
        RECT 0.000 0.000 9.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.600 3.950 0.850 7.250 ;
        RECT 3.150 5.800 3.400 7.250 ;
        RECT 1.150 5.550 3.400 5.800 ;
        RECT 5.700 5.600 5.950 7.250 ;
        RECT 1.150 4.550 1.400 5.550 ;
        RECT 5.700 5.350 6.200 5.600 ;
        RECT 2.600 4.800 3.100 5.100 ;
        RECT 1.100 4.250 1.550 4.550 ;
        RECT 1.850 4.250 2.350 4.550 ;
        RECT 0.500 3.900 0.850 3.950 ;
        RECT 0.350 3.600 0.850 3.900 ;
        RECT 0.450 3.550 0.850 3.600 ;
        RECT 0.600 1.050 0.850 3.550 ;
        RECT 1.150 2.400 1.400 4.250 ;
        RECT 2.700 2.950 3.000 4.800 ;
        RECT 3.450 4.250 3.950 4.550 ;
        RECT 5.200 4.250 5.700 4.550 ;
        RECT 4.500 3.600 5.000 3.900 ;
        RECT 5.950 2.950 6.200 5.350 ;
        RECT 6.450 5.400 6.700 7.250 ;
        RECT 6.450 5.200 6.850 5.400 ;
        RECT 8.150 5.250 8.400 7.250 ;
        RECT 8.150 5.200 8.550 5.250 ;
        RECT 6.450 5.150 6.950 5.200 ;
        RECT 6.450 4.900 7.800 5.150 ;
        RECT 6.450 4.850 6.850 4.900 ;
        RECT 6.750 3.600 7.250 3.900 ;
        RECT 2.700 2.650 6.200 2.950 ;
        RECT 1.150 2.150 3.400 2.400 ;
        RECT 5.950 2.300 6.200 2.650 ;
        RECT 7.500 2.400 7.800 4.900 ;
        RECT 3.150 1.050 3.400 2.150 ;
        RECT 5.700 2.050 6.200 2.300 ;
        RECT 6.450 2.150 7.800 2.400 ;
        RECT 8.150 4.900 8.650 5.200 ;
        RECT 8.150 4.850 8.550 4.900 ;
        RECT 5.700 1.050 5.950 2.050 ;
        RECT 6.450 1.050 6.700 2.150 ;
        RECT 8.150 1.050 8.400 4.850 ;
      LAYER Via1 ;
        RECT 1.950 4.250 2.250 4.550 ;
        RECT 0.450 3.600 0.750 3.900 ;
        RECT 3.550 4.250 3.850 4.550 ;
        RECT 5.300 4.250 5.600 4.550 ;
        RECT 4.600 3.600 4.900 3.900 ;
        RECT 6.550 4.900 6.850 5.200 ;
        RECT 6.850 3.600 7.150 3.900 ;
        RECT 8.250 4.900 8.550 5.200 ;
      LAYER Metal2 ;
        RECT 6.500 5.200 6.900 5.250 ;
        RECT 6.450 4.900 6.950 5.200 ;
        RECT 6.500 4.850 6.900 4.900 ;
        RECT 0.350 3.900 0.850 3.950 ;
        RECT 4.550 3.900 4.950 3.950 ;
        RECT 6.750 3.900 7.250 3.950 ;
        RECT 0.350 3.600 7.250 3.900 ;
        RECT 0.350 3.550 0.850 3.600 ;
        RECT 4.550 3.550 4.950 3.600 ;
        RECT 6.750 3.550 7.250 3.600 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dlat_1


MACRO gf180mcu_osu_sc_gp12t3v3__tbuf_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tbuf_1 ;
  SIZE 5.200 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN EN
    ANTENNAGATEAREA 1.020000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.000 2.300 3.500 2.700 ;
    END
  END EN
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.450 3.550 2.950 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.135000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 5.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 5.200 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.550 5.550 3.800 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.242500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.550 0.700 3.800 1.900 ;
        RECT 0.000 0.000 5.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.750 0.800 7.250 ;
        RECT 2.800 5.800 3.050 7.250 ;
        RECT 1.950 5.550 3.050 5.800 ;
        RECT 1.950 4.600 2.200 5.550 ;
        RECT 4.400 5.200 4.650 7.250 ;
        RECT 2.450 4.900 2.950 5.200 ;
        RECT 4.300 4.900 4.800 5.200 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.950 4.350 2.800 4.600 ;
        RECT 2.550 3.900 2.800 4.350 ;
        RECT 0.550 3.450 2.000 3.750 ;
        RECT 2.450 3.600 2.950 3.900 ;
        RECT 0.550 1.050 0.800 3.450 ;
        RECT 2.550 3.100 2.800 3.600 ;
        RECT 1.950 2.850 2.800 3.100 ;
        RECT 1.950 1.900 2.200 2.850 ;
        RECT 3.000 2.350 3.500 2.650 ;
        RECT 1.950 1.650 3.050 1.900 ;
        RECT 2.800 1.050 3.050 1.650 ;
        RECT 4.400 1.050 4.650 4.900 ;
      LAYER Via1 ;
        RECT 2.550 4.900 2.850 5.200 ;
        RECT 4.400 4.900 4.700 5.200 ;
        RECT 1.150 4.250 1.450 4.550 ;
        RECT 2.550 3.600 2.850 3.900 ;
        RECT 3.100 2.350 3.400 2.650 ;
      LAYER Metal2 ;
        RECT 2.450 5.200 2.950 5.250 ;
        RECT 4.300 5.200 4.800 5.250 ;
        RECT 2.450 4.900 4.800 5.200 ;
        RECT 2.450 4.850 2.950 4.900 ;
        RECT 4.300 4.850 4.800 4.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tbuf_1


MACRO gf180mcu_osu_sc_gp12t3v3__inv_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_2 ;
  SIZE 3.200 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.650 3.550 1.150 3.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 1.500 4.200 2.000 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.460000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.200 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.300 5.550 2.550 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 0.000 0.000 3.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.650 1.650 7.250 ;
        RECT 1.400 4.550 1.850 4.650 ;
        RECT 1.400 4.250 2.000 4.550 ;
        RECT 1.400 4.100 1.850 4.250 ;
        RECT 0.650 3.600 1.150 3.900 ;
        RECT 1.400 1.050 1.650 4.100 ;
      LAYER Via1 ;
        RECT 1.600 4.250 1.900 4.550 ;
        RECT 0.750 3.600 1.050 3.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__inv_2


MACRO gf180mcu_osu_sc_gp12t3v3__aoi21_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi21_1 ;
  SIZE 3.900 BY 8.300 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 3.550 1.100 3.950 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.600 4.200 2.100 4.600 ;
    END
  END A1
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.350 3.550 2.850 3.950 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.317500 ;
    PORT
      LAYER Metal2 ;
        RECT 3.000 4.850 3.500 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.947500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.900 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.900 8.300 ;
        RECT 1.400 6.300 1.650 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.862500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 0.700 0.950 1.900 ;
        RECT 2.950 0.700 3.200 1.900 ;
        RECT 0.000 0.000 3.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 6.050 0.800 7.250 ;
        RECT 2.250 6.050 2.500 7.250 ;
        RECT 0.550 5.800 2.500 6.050 ;
        RECT 3.100 5.200 3.350 7.250 ;
        RECT 3.000 4.900 3.500 5.200 ;
        RECT 1.600 4.250 2.100 4.550 ;
        RECT 0.600 3.600 1.100 3.900 ;
        RECT 2.350 3.600 2.850 3.900 ;
        RECT 3.100 2.900 3.350 4.900 ;
        RECT 2.100 2.650 3.350 2.900 ;
        RECT 2.100 1.050 2.350 2.650 ;
      LAYER Via1 ;
        RECT 3.100 4.900 3.400 5.200 ;
        RECT 1.700 4.250 2.000 4.550 ;
        RECT 0.700 3.600 1.000 3.900 ;
        RECT 2.450 3.600 2.750 3.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi21_1


MACRO gf180mcu_osu_sc_gp12t3v3__buf_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_1 ;
  SIZE 3.100 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.150 4.850 2.650 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.610000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.100 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.100 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.142500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 0.000 0.000 3.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.200 2.500 7.250 ;
        RECT 2.150 4.900 2.650 5.200 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 1.050 2.500 4.900 ;
      LAYER Via1 ;
        RECT 2.250 4.900 2.550 5.200 ;
        RECT 1.150 4.250 1.450 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_1


MACRO gf180mcu_osu_sc_gp12t3v3__dff_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dff_1 ;
  SIZE 13.000 BY 8.300 ;
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.900 3.900 2.400 3.950 ;
        RECT 1.750 3.600 2.550 3.900 ;
        RECT 1.900 3.550 2.400 3.600 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.250 4.550 3.700 4.600 ;
        RECT 6.050 4.550 6.550 4.600 ;
        RECT 7.700 4.550 8.100 4.600 ;
        RECT 3.250 4.250 8.150 4.550 ;
        RECT 3.250 4.200 3.700 4.250 ;
        RECT 6.050 4.200 6.550 4.250 ;
        RECT 7.700 4.200 8.100 4.250 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.200 5.200 12.600 5.250 ;
        RECT 12.150 4.900 12.650 5.200 ;
        RECT 12.200 4.850 12.600 4.900 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 0.765000 ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.450 4.550 11.850 4.600 ;
        RECT 11.400 4.250 11.900 4.550 ;
        RECT 11.450 4.200 11.850 4.250 ;
    END
  END QN
  PIN VDD
    ANTENNADIFFAREA 7.965001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 13.000 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 13.000 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 4.450 5.550 4.700 7.600 ;
        RECT 7.250 6.300 7.500 7.600 ;
        RECT 8.850 5.550 9.100 7.600 ;
        RECT 11.300 5.550 11.550 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 5.595000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 4.450 0.700 4.700 1.500 ;
        RECT 7.250 0.700 7.500 1.900 ;
        RECT 8.850 0.700 9.100 1.550 ;
        RECT 11.300 0.700 11.550 1.900 ;
        RECT 0.000 0.000 13.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.700 0.800 7.250 ;
        RECT 3.050 5.300 3.300 7.250 ;
        RECT 5.850 6.300 6.100 7.250 ;
        RECT 1.400 5.050 3.300 5.300 ;
        RECT 4.950 6.050 6.100 6.300 ;
        RECT 1.400 4.550 1.650 5.050 ;
        RECT 4.050 4.900 4.550 5.200 ;
        RECT 1.050 4.250 1.650 4.550 ;
        RECT 2.600 4.250 3.750 4.550 ;
        RECT 0.500 2.200 0.800 2.700 ;
        RECT 1.400 2.600 1.650 4.250 ;
        RECT 3.350 4.200 3.650 4.250 ;
        RECT 1.900 3.600 2.400 3.900 ;
        RECT 2.900 2.950 3.400 3.250 ;
        RECT 4.150 2.600 4.450 4.900 ;
        RECT 4.950 3.800 5.200 6.050 ;
        RECT 6.700 4.900 7.200 5.200 ;
        RECT 8.100 5.100 8.350 7.250 ;
        RECT 4.900 3.550 5.200 3.800 ;
        RECT 5.500 4.250 6.550 4.550 ;
        RECT 1.400 2.350 2.400 2.600 ;
        RECT 0.550 1.050 0.800 2.200 ;
        RECT 2.000 1.900 2.400 2.350 ;
        RECT 4.050 2.300 4.550 2.600 ;
        RECT 4.900 1.950 5.150 3.550 ;
        RECT 5.500 2.650 5.800 4.250 ;
        RECT 6.800 3.900 7.100 4.900 ;
        RECT 8.100 4.850 8.900 5.100 ;
        RECT 7.650 4.250 8.150 4.550 ;
        RECT 8.600 3.900 8.900 4.850 ;
        RECT 6.750 3.600 7.300 3.900 ;
        RECT 8.100 3.650 8.900 3.900 ;
        RECT 6.800 3.550 7.200 3.600 ;
        RECT 8.100 2.850 8.400 3.650 ;
        RECT 9.050 3.250 9.350 3.350 ;
        RECT 9.700 3.250 9.950 7.250 ;
        RECT 10.450 4.550 10.700 7.250 ;
        RECT 12.150 5.250 12.400 7.250 ;
        RECT 12.150 4.900 12.650 5.250 ;
        RECT 12.150 4.850 12.600 4.900 ;
        RECT 10.450 4.250 11.900 4.550 ;
        RECT 8.950 2.950 9.450 3.250 ;
        RECT 9.700 2.950 11.150 3.250 ;
        RECT 5.400 2.250 5.900 2.650 ;
        RECT 2.000 1.650 3.300 1.900 ;
        RECT 4.900 1.700 6.250 1.950 ;
        RECT 3.050 1.050 3.300 1.650 ;
        RECT 5.850 1.650 6.250 1.700 ;
        RECT 5.850 1.050 6.100 1.650 ;
        RECT 8.100 1.050 8.350 2.850 ;
        RECT 9.050 2.100 9.350 2.950 ;
        RECT 8.950 1.800 9.450 2.100 ;
        RECT 9.700 1.050 9.950 2.950 ;
        RECT 11.550 2.400 11.800 4.250 ;
        RECT 10.450 2.150 11.800 2.400 ;
        RECT 10.450 1.050 10.700 2.150 ;
        RECT 12.150 1.050 12.400 4.850 ;
      LAYER Via1 ;
        RECT 3.350 4.250 3.650 4.550 ;
        RECT 0.500 2.300 0.800 2.600 ;
        RECT 2.000 3.600 2.300 3.900 ;
        RECT 3.000 2.950 3.300 3.250 ;
        RECT 6.800 4.900 7.100 5.200 ;
        RECT 6.150 4.250 6.450 4.550 ;
        RECT 4.150 2.300 4.450 2.600 ;
        RECT 7.750 4.250 8.050 4.550 ;
        RECT 6.850 3.600 7.150 3.900 ;
        RECT 12.250 4.900 12.550 5.200 ;
        RECT 11.500 4.250 11.800 4.550 ;
        RECT 8.100 2.950 8.400 3.250 ;
        RECT 10.750 2.950 11.050 3.250 ;
        RECT 9.050 1.800 9.350 2.100 ;
      LAYER Metal2 ;
        RECT 6.750 5.200 7.150 5.250 ;
        RECT 6.700 4.900 9.900 5.200 ;
        RECT 6.750 4.850 7.150 4.900 ;
        RECT 6.800 3.900 7.200 3.950 ;
        RECT 6.750 3.600 7.250 3.900 ;
        RECT 6.800 3.550 7.200 3.600 ;
        RECT 2.950 3.250 3.350 3.300 ;
        RECT 8.050 3.250 8.450 3.300 ;
        RECT 9.600 3.250 9.900 4.900 ;
        RECT 10.700 3.250 11.100 3.300 ;
        RECT 2.900 2.950 8.550 3.250 ;
        RECT 9.600 2.950 11.150 3.250 ;
        RECT 2.950 2.900 3.350 2.950 ;
        RECT 8.050 2.900 8.450 2.950 ;
        RECT 10.700 2.900 11.100 2.950 ;
        RECT 0.450 2.600 0.850 2.650 ;
        RECT 4.100 2.600 4.500 2.650 ;
        RECT 0.400 2.300 4.550 2.600 ;
        RECT 0.450 2.250 0.850 2.300 ;
        RECT 4.100 2.250 4.500 2.300 ;
        RECT 9.000 2.100 9.400 2.150 ;
        RECT 5.800 1.950 6.200 2.000 ;
        RECT 8.500 1.950 9.450 2.100 ;
        RECT 5.750 1.800 9.450 1.950 ;
        RECT 5.750 1.750 9.400 1.800 ;
        RECT 5.750 1.650 8.800 1.750 ;
        RECT 5.800 1.600 6.200 1.650 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dff_1


MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_4 ;
  SIZE 5.600 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.805000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.850 5.250 4.350 5.300 ;
        RECT 3.800 4.950 4.350 5.250 ;
        RECT 3.850 4.900 4.350 4.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 4.070000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 5.600 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 5.600 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
        RECT 4.800 5.550 5.050 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.710000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 0.000 0.000 5.600 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.250 2.500 7.250 ;
        RECT 3.950 5.250 4.200 7.250 ;
        RECT 2.250 4.950 4.350 5.250 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 2.400 2.500 4.950 ;
        RECT 3.950 2.400 4.200 4.950 ;
        RECT 2.250 2.150 4.200 2.400 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
      LAYER Via1 ;
        RECT 3.950 4.950 4.250 5.250 ;
        RECT 1.150 4.250 1.450 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_4


MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_2 ;
  SIZE 3.200 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.650 3.550 1.150 3.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 1.500 4.450 2.000 4.850 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.122500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.200 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.300 5.550 2.550 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 0.000 0.000 3.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.900 1.650 7.250 ;
        RECT 1.400 4.800 1.850 4.900 ;
        RECT 1.400 4.500 2.000 4.800 ;
        RECT 1.400 4.350 1.850 4.500 ;
        RECT 0.650 3.600 1.150 3.900 ;
        RECT 1.400 1.050 1.650 4.350 ;
      LAYER Via1 ;
        RECT 1.600 4.500 1.900 4.800 ;
        RECT 0.750 3.600 1.050 3.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkinv_2


MACRO gf180mcu_osu_sc_gp12t3v3__inv_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_1 ;
  SIZE 2.200 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.550 4.850 1.050 5.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 3.550 1.800 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 2.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 2.200 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.762500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.900 1.050 5.200 ;
        RECT 1.400 3.900 1.650 7.250 ;
        RECT 1.300 3.600 1.800 3.900 ;
        RECT 1.400 1.050 1.650 3.600 ;
      LAYER Via1 ;
        RECT 0.650 4.900 0.950 5.200 ;
        RECT 1.400 3.600 1.700 3.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__inv_1


MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_1 ;
  SIZE 3.100 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.150 4.850 2.650 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.610000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.100 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.100 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.142500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 0.000 0.000 3.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.200 2.500 7.250 ;
        RECT 2.150 4.900 2.650 5.200 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 1.050 2.500 4.900 ;
      LAYER Via1 ;
        RECT 2.250 4.900 2.550 5.200 ;
        RECT 1.150 4.250 1.450 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_1


MACRO gf180mcu_osu_sc_gp12t3v3__buf_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_8 ;
  SIZE 9.000 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 5.610001 ;
    PORT
      LAYER Metal2 ;
        RECT 7.200 4.950 7.750 5.250 ;
        RECT 7.250 4.850 7.750 4.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 6.615000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 9.000 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 9.000 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
        RECT 4.800 5.550 5.050 7.600 ;
        RECT 6.500 5.550 6.750 7.600 ;
        RECT 8.200 5.550 8.450 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.900 ;
        RECT 8.200 0.700 8.450 1.900 ;
        RECT 0.000 0.000 9.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.250 2.500 7.250 ;
        RECT 3.950 5.250 4.200 7.250 ;
        RECT 5.650 5.250 5.900 7.250 ;
        RECT 7.350 5.250 7.600 7.250 ;
        RECT 2.250 5.200 7.600 5.250 ;
        RECT 2.250 4.950 7.750 5.200 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 2.400 2.500 4.950 ;
        RECT 3.950 2.400 4.200 4.950 ;
        RECT 5.650 2.400 5.900 4.950 ;
        RECT 7.250 4.900 7.750 4.950 ;
        RECT 7.350 2.400 7.600 4.900 ;
        RECT 2.250 2.150 7.600 2.400 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
        RECT 5.650 1.050 5.900 2.150 ;
        RECT 7.350 1.050 7.600 2.150 ;
      LAYER Via1 ;
        RECT 1.150 4.250 1.450 4.550 ;
        RECT 7.350 4.900 7.650 5.200 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_8


MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_16 ;
  SIZE 15.800 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 11.220001 ;
    PORT
      LAYER Metal2 ;
        RECT 14.050 5.250 14.550 5.300 ;
        RECT 14.000 4.950 14.550 5.250 ;
        RECT 14.050 4.900 14.550 4.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 12.380001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 15.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 15.800 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
        RECT 4.800 5.550 5.050 7.600 ;
        RECT 6.500 5.550 6.750 7.600 ;
        RECT 8.200 5.550 8.450 7.600 ;
        RECT 9.900 5.550 10.150 7.600 ;
        RECT 11.600 5.550 11.850 7.600 ;
        RECT 13.300 5.550 13.550 7.600 ;
        RECT 15.000 5.550 15.250 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.215000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.900 ;
        RECT 8.200 0.700 8.450 1.900 ;
        RECT 9.900 0.700 10.150 1.900 ;
        RECT 11.600 0.700 11.850 1.900 ;
        RECT 13.300 0.700 13.550 1.900 ;
        RECT 15.000 0.700 15.250 1.900 ;
        RECT 0.000 0.000 15.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.250 2.500 7.250 ;
        RECT 3.950 5.250 4.200 7.250 ;
        RECT 5.650 5.250 5.900 7.250 ;
        RECT 7.350 5.250 7.600 7.250 ;
        RECT 9.050 5.250 9.300 7.250 ;
        RECT 10.750 5.250 11.000 7.250 ;
        RECT 12.450 5.250 12.700 7.250 ;
        RECT 14.150 5.250 14.400 7.250 ;
        RECT 2.250 4.950 14.550 5.250 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 2.400 2.500 4.950 ;
        RECT 3.950 2.400 4.200 4.950 ;
        RECT 5.650 2.400 5.900 4.950 ;
        RECT 7.350 2.400 7.600 4.950 ;
        RECT 9.050 2.400 9.300 4.950 ;
        RECT 10.750 2.400 11.000 4.950 ;
        RECT 12.450 2.400 12.700 4.950 ;
        RECT 14.150 2.400 14.400 4.950 ;
        RECT 2.250 2.150 14.400 2.400 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
        RECT 5.650 1.050 5.900 2.150 ;
        RECT 7.350 1.050 7.600 2.150 ;
        RECT 9.050 1.050 9.300 2.150 ;
        RECT 10.750 1.050 11.000 2.150 ;
        RECT 12.450 1.050 12.700 2.150 ;
        RECT 14.150 1.050 14.400 2.150 ;
      LAYER Via1 ;
        RECT 14.150 4.950 14.450 5.250 ;
        RECT 1.150 4.250 1.450 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_16


MACRO gf180mcu_osu_sc_gp12t3v3__dlatn_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dlatn_1 ;
  SIZE 10.700 BY 8.300 ;
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.850 4.200 2.350 4.600 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.050 2.600 7.550 3.000 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.900 5.200 10.300 5.250 ;
        RECT 9.850 4.900 10.350 5.200 ;
        RECT 9.900 4.850 10.300 4.900 ;
    END
  END Q
  PIN VDD
    ANTENNADIFFAREA 6.355000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 10.700 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 10.700 8.300 ;
        RECT 1.450 6.350 1.700 7.600 ;
        RECT 4.850 5.550 5.100 7.600 ;
        RECT 7.400 5.550 7.650 7.600 ;
        RECT 9.000 5.550 9.250 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.782500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 0.700 1.850 1.900 ;
        RECT 4.700 0.700 5.100 1.900 ;
        RECT 7.400 0.700 7.650 1.900 ;
        RECT 9.000 0.700 9.250 1.900 ;
        RECT 0.000 0.000 10.700 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.600 3.950 0.850 7.250 ;
        RECT 3.150 5.800 3.400 7.250 ;
        RECT 1.150 5.550 3.400 5.800 ;
        RECT 5.700 5.600 5.950 7.250 ;
        RECT 1.150 4.550 1.400 5.550 ;
        RECT 5.700 5.350 6.200 5.600 ;
        RECT 2.600 4.800 3.100 5.100 ;
        RECT 1.100 4.250 1.550 4.550 ;
        RECT 1.850 4.250 2.350 4.550 ;
        RECT 0.500 3.900 0.850 3.950 ;
        RECT 0.350 3.600 0.850 3.900 ;
        RECT 0.450 3.550 0.850 3.600 ;
        RECT 0.600 1.050 0.850 3.550 ;
        RECT 1.150 2.400 1.400 4.250 ;
        RECT 2.700 2.950 3.000 4.800 ;
        RECT 3.450 4.250 3.950 4.550 ;
        RECT 5.200 4.250 5.700 4.550 ;
        RECT 4.500 3.600 5.000 3.900 ;
        RECT 5.950 2.950 6.200 5.350 ;
        RECT 6.550 4.600 6.800 7.250 ;
        RECT 8.150 5.400 8.400 7.250 ;
        RECT 8.150 5.200 8.550 5.400 ;
        RECT 9.850 5.250 10.100 7.250 ;
        RECT 9.850 5.200 10.250 5.250 ;
        RECT 8.150 5.150 8.650 5.200 ;
        RECT 8.150 4.900 9.500 5.150 ;
        RECT 8.150 4.850 8.550 4.900 ;
        RECT 6.550 4.550 6.950 4.600 ;
        RECT 6.450 4.250 6.950 4.550 ;
        RECT 2.700 2.650 6.200 2.950 ;
        RECT 1.150 2.150 3.400 2.400 ;
        RECT 5.950 2.300 6.200 2.650 ;
        RECT 3.150 1.050 3.400 2.150 ;
        RECT 5.700 2.050 6.200 2.300 ;
        RECT 6.550 4.200 6.950 4.250 ;
        RECT 5.700 1.050 5.950 2.050 ;
        RECT 6.550 1.050 6.800 4.200 ;
        RECT 8.450 3.600 8.950 3.900 ;
        RECT 7.050 2.650 7.550 2.950 ;
        RECT 9.200 2.400 9.500 4.900 ;
        RECT 8.150 2.150 9.500 2.400 ;
        RECT 9.850 4.900 10.350 5.200 ;
        RECT 9.850 4.850 10.250 4.900 ;
        RECT 8.150 1.050 8.400 2.150 ;
        RECT 9.850 1.050 10.100 4.850 ;
      LAYER Via1 ;
        RECT 1.950 4.250 2.250 4.550 ;
        RECT 0.450 3.600 0.750 3.900 ;
        RECT 3.550 4.250 3.850 4.550 ;
        RECT 5.300 4.250 5.600 4.550 ;
        RECT 4.600 3.600 4.900 3.900 ;
        RECT 8.250 4.900 8.550 5.200 ;
        RECT 6.550 4.250 6.850 4.550 ;
        RECT 8.550 3.600 8.850 3.900 ;
        RECT 7.150 2.650 7.450 2.950 ;
        RECT 9.950 4.900 10.250 5.200 ;
      LAYER Metal2 ;
        RECT 8.200 5.200 8.600 5.250 ;
        RECT 8.150 4.900 8.650 5.200 ;
        RECT 8.200 4.850 8.600 4.900 ;
        RECT 3.500 4.550 3.900 4.600 ;
        RECT 5.200 4.550 5.700 4.600 ;
        RECT 6.450 4.550 6.950 4.600 ;
        RECT 3.450 4.250 6.950 4.550 ;
        RECT 3.500 4.200 3.900 4.250 ;
        RECT 5.200 4.200 5.700 4.250 ;
        RECT 6.450 4.200 6.950 4.250 ;
        RECT 0.350 3.900 0.850 3.950 ;
        RECT 4.550 3.900 4.950 3.950 ;
        RECT 8.450 3.900 8.950 3.950 ;
        RECT 0.350 3.600 8.950 3.900 ;
        RECT 0.350 3.550 0.850 3.600 ;
        RECT 4.550 3.550 4.950 3.600 ;
        RECT 8.450 3.550 8.950 3.600 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dlatn_1


MACRO gf180mcu_osu_sc_gp12t3v3__xor2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__xor2_1 ;
  SIZE 6.200 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 2.600 1.700 2.650 ;
        RECT 1.250 2.300 1.750 2.600 ;
        RECT 1.300 2.250 1.700 2.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.000 3.900 2.400 3.950 ;
        RECT 4.650 3.900 5.050 3.950 ;
        RECT 1.950 3.600 2.450 3.900 ;
        RECT 4.600 3.600 5.100 3.900 ;
        RECT 2.000 3.550 2.400 3.600 ;
        RECT 4.650 3.550 5.050 3.600 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 2.192500 ;
    PORT
      LAYER Metal2 ;
        RECT 2.900 5.900 3.200 6.050 ;
        RECT 2.850 5.500 3.250 5.900 ;
        RECT 2.900 2.000 3.200 5.500 ;
        RECT 2.800 1.600 3.300 2.000 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.557500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 6.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 6.200 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 4.500 5.550 4.750 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.622500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 4.500 0.700 4.750 1.900 ;
        RECT 0.000 0.000 6.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.550 0.800 7.250 ;
        RECT 2.950 5.950 3.200 7.250 ;
        RECT 2.900 5.450 3.200 5.950 ;
        RECT 5.350 5.200 5.600 7.250 ;
        RECT 2.550 4.900 5.600 5.200 ;
        RECT 0.550 4.250 4.050 4.550 ;
        RECT 0.550 1.050 0.800 4.250 ;
        RECT 1.950 3.600 5.100 3.900 ;
        RECT 5.350 2.600 5.600 4.900 ;
        RECT 1.250 2.300 1.750 2.600 ;
        RECT 4.050 2.300 5.600 2.600 ;
        RECT 2.900 1.500 3.200 2.050 ;
        RECT 2.950 1.050 3.200 1.500 ;
        RECT 5.350 1.050 5.600 2.300 ;
      LAYER Via1 ;
        RECT 2.900 5.550 3.200 5.850 ;
        RECT 2.050 3.600 2.350 3.900 ;
        RECT 4.700 3.600 5.000 3.900 ;
        RECT 1.350 2.300 1.650 2.600 ;
        RECT 2.900 1.650 3.200 1.950 ;
  END
END gf180mcu_osu_sc_gp12t3v3__xor2_1


MACRO gf180mcu_osu_sc_gp12t3v3__fill_4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_4 ;
  SIZE 0.900 BY 8.300 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.600 0.400 8.300 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 0.400 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 5.100 0.400 8.300 ;
  END
END gf180mcu_osu_sc_gp12t3v3__fill_4


MACRO gf180mcu_osu_sc_gp12t3v3__tinv_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tinv_1 ;
  SIZE 3.650 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.450 4.850 1.950 5.250 ;
    END
  END A
  PIN EN
    ANTENNAGATEAREA 1.020000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.000 2.600 1.500 2.650 ;
        RECT 2.700 2.600 3.200 2.650 ;
        RECT 1.000 2.300 3.200 2.600 ;
        RECT 1.000 2.250 1.500 2.300 ;
        RECT 2.700 2.250 3.200 2.300 ;
    END
  END EN
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.050 3.550 2.550 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.947500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.650 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.650 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.480000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 0.000 0.000 3.650 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 5.800 0.800 7.250 ;
        RECT 2.800 5.800 3.050 7.250 ;
        RECT 0.500 5.550 0.800 5.800 ;
        RECT 2.200 5.550 3.050 5.800 ;
        RECT 0.500 4.550 0.750 5.550 ;
        RECT 1.450 4.900 1.950 5.200 ;
        RECT 0.350 4.250 0.850 4.550 ;
        RECT 0.500 2.150 0.750 4.250 ;
        RECT 2.200 3.900 2.450 5.550 ;
        RECT 2.700 4.900 3.200 5.200 ;
        RECT 2.050 3.600 2.600 3.900 ;
        RECT 1.000 2.300 1.500 2.600 ;
        RECT 0.500 1.900 0.800 2.150 ;
        RECT 0.550 1.050 0.800 1.900 ;
        RECT 2.200 1.900 2.450 3.600 ;
        RECT 2.700 2.300 3.200 2.600 ;
        RECT 2.200 1.650 3.050 1.900 ;
        RECT 2.800 1.050 3.050 1.650 ;
      LAYER Via1 ;
        RECT 1.550 4.900 1.850 5.200 ;
        RECT 0.450 4.250 0.750 4.550 ;
        RECT 2.800 4.900 3.100 5.200 ;
        RECT 2.150 3.600 2.450 3.900 ;
        RECT 1.100 2.300 1.400 2.600 ;
        RECT 2.800 2.300 3.100 2.600 ;
      LAYER Metal2 ;
        RECT 2.700 4.850 3.200 5.250 ;
        RECT 0.350 4.550 0.850 4.600 ;
        RECT 2.800 4.550 3.100 4.850 ;
        RECT 0.350 4.250 3.100 4.550 ;
        RECT 0.350 4.200 0.850 4.250 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tinv_1


MACRO gf180mcu_osu_sc_gp12t3v3__fill_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_1 ;
  SIZE 0.900 BY 8.300 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.600 0.100 8.300 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 0.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 5.100 0.100 8.300 ;
  END
END gf180mcu_osu_sc_gp12t3v3__fill_1


MACRO gf180mcu_osu_sc_gp12t3v3__oai31_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai31_1 ;
  SIZE 4.800 BY 8.300 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.950 2.900 1.450 3.300 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.800 2.900 2.300 3.300 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.550 4.200 3.050 4.600 ;
    END
  END A2
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.100 2.900 3.600 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.360000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.750 4.850 4.250 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.050000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 4.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 4.800 8.300 ;
        RECT 1.050 5.550 1.300 7.600 ;
        RECT 3.850 5.550 4.100 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.242500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.600 ;
        RECT 0.000 0.000 4.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.000 5.200 3.250 7.250 ;
        RECT 3.000 4.900 4.250 5.200 ;
        RECT 2.550 4.250 3.050 4.550 ;
        RECT 0.950 2.950 1.450 3.250 ;
        RECT 1.800 2.950 2.300 3.250 ;
        RECT 3.100 2.950 3.600 3.250 ;
        RECT 3.850 2.600 4.100 4.900 ;
        RECT 3.850 2.350 4.200 2.600 ;
        RECT 1.400 1.850 3.350 2.100 ;
        RECT 1.400 1.050 1.650 1.850 ;
        RECT 3.100 1.050 3.350 1.850 ;
        RECT 3.950 1.050 4.200 2.350 ;
      LAYER Via1 ;
        RECT 3.850 4.900 4.150 5.200 ;
        RECT 2.650 4.250 2.950 4.550 ;
        RECT 1.050 2.950 1.350 3.250 ;
        RECT 1.900 2.950 2.200 3.250 ;
        RECT 3.200 2.950 3.500 3.250 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai31_1


MACRO gf180mcu_osu_sc_gp12t3v3__buf_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_16 ;
  SIZE 15.800 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 11.220001 ;
    PORT
      LAYER Metal2 ;
        RECT 14.000 4.950 14.550 5.250 ;
        RECT 14.050 4.850 14.550 4.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 12.380001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 15.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 15.800 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
        RECT 4.800 5.550 5.050 7.600 ;
        RECT 6.500 5.550 6.750 7.600 ;
        RECT 8.200 5.550 8.450 7.600 ;
        RECT 9.900 5.550 10.150 7.600 ;
        RECT 11.600 5.550 11.850 7.600 ;
        RECT 13.300 5.550 13.550 7.600 ;
        RECT 15.000 5.550 15.250 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.215000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.900 ;
        RECT 8.200 0.700 8.450 1.900 ;
        RECT 9.900 0.700 10.150 1.900 ;
        RECT 11.600 0.700 11.850 1.900 ;
        RECT 13.300 0.700 13.550 1.900 ;
        RECT 15.000 0.700 15.250 1.900 ;
        RECT 0.000 0.000 15.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.250 2.500 7.250 ;
        RECT 3.950 5.250 4.200 7.250 ;
        RECT 5.650 5.250 5.900 7.250 ;
        RECT 7.350 5.250 7.600 7.250 ;
        RECT 9.050 5.250 9.300 7.250 ;
        RECT 10.750 5.250 11.000 7.250 ;
        RECT 12.450 5.250 12.700 7.250 ;
        RECT 14.150 5.250 14.400 7.250 ;
        RECT 2.250 5.200 14.400 5.250 ;
        RECT 2.250 4.950 14.550 5.200 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 2.400 2.500 4.950 ;
        RECT 3.950 2.400 4.200 4.950 ;
        RECT 5.650 2.400 5.900 4.950 ;
        RECT 7.350 2.400 7.600 4.950 ;
        RECT 9.050 2.400 9.300 4.950 ;
        RECT 10.750 2.400 11.000 4.950 ;
        RECT 12.450 2.400 12.700 4.950 ;
        RECT 14.050 4.900 14.550 4.950 ;
        RECT 14.150 2.400 14.400 4.900 ;
        RECT 2.250 2.150 14.400 2.400 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
        RECT 5.650 1.050 5.900 2.150 ;
        RECT 7.350 1.050 7.600 2.150 ;
        RECT 9.050 1.050 9.300 2.150 ;
        RECT 10.750 1.050 11.000 2.150 ;
        RECT 12.450 1.050 12.700 2.150 ;
        RECT 14.150 1.050 14.400 2.150 ;
      LAYER Via1 ;
        RECT 1.150 4.250 1.450 4.550 ;
        RECT 14.150 4.900 14.450 5.200 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_16


MACRO gf180mcu_osu_sc_gp12t3v3__buf_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_2 ;
  SIZE 3.900 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 2.150 4.850 2.650 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.460000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.900 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.900 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.567500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 0.000 0.000 3.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.200 2.500 7.250 ;
        RECT 2.150 4.900 2.650 5.200 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 1.050 2.500 4.900 ;
      LAYER Via1 ;
        RECT 2.250 4.900 2.550 5.200 ;
        RECT 1.150 4.250 1.450 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_2


MACRO gf180mcu_osu_sc_gp12t3v3__mux2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__mux2_1 ;
  SIZE 4.800 BY 8.300 ;
  PIN A
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.350 3.550 2.850 3.950 ;
    END
  END A
  PIN B
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.750 4.200 4.250 4.600 ;
    END
  END B
  PIN Sel
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.550 2.900 1.050 3.300 ;
    END
  END Sel
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 3.000 4.850 3.500 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.862500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 4.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 4.800 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.437500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 4.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.550 1.650 7.250 ;
        RECT 1.400 4.250 2.000 4.550 ;
        RECT 0.550 2.950 1.050 3.250 ;
        RECT 1.400 2.600 1.650 4.250 ;
        RECT 2.250 3.950 2.500 7.250 ;
        RECT 3.100 5.250 3.350 7.250 ;
        RECT 3.000 4.850 3.500 5.250 ;
        RECT 2.250 3.550 2.850 3.950 ;
        RECT 1.400 2.300 2.000 2.600 ;
        RECT 1.400 1.050 1.650 2.300 ;
        RECT 2.250 1.050 2.500 3.550 ;
        RECT 3.100 1.050 3.350 4.850 ;
        RECT 3.950 4.600 4.200 7.250 ;
        RECT 3.750 4.200 4.250 4.600 ;
        RECT 3.950 1.050 4.200 4.200 ;
      LAYER Via1 ;
        RECT 0.650 2.950 0.950 3.250 ;
        RECT 3.100 4.900 3.400 5.200 ;
        RECT 2.450 3.600 2.750 3.900 ;
        RECT 3.850 4.250 4.150 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__mux2_1


MACRO gf180mcu_osu_sc_gp12t3v3__nand2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nand2_1 ;
  SIZE 3.100 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 3.550 1.100 3.950 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.900 2.900 2.400 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.360000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 4.200 1.800 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.375000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.100 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.100 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.100000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.700 2.350 1.900 ;
        RECT 0.000 0.000 3.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.550 1.650 7.250 ;
        RECT 1.300 4.250 1.800 4.550 ;
        RECT 0.600 3.600 1.100 3.900 ;
        RECT 1.400 2.250 1.650 4.250 ;
        RECT 1.900 2.950 2.400 3.250 ;
        RECT 0.700 2.000 1.650 2.250 ;
        RECT 0.700 1.050 0.950 2.000 ;
      LAYER Via1 ;
        RECT 1.400 4.250 1.700 4.550 ;
        RECT 0.700 3.600 1.000 3.900 ;
        RECT 2.000 2.950 2.300 3.250 ;
  END
END gf180mcu_osu_sc_gp12t3v3__nand2_1


MACRO gf180mcu_osu_sc_gp12t3v3__oai21_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai21_1 ;
  SIZE 3.900 BY 8.300 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.450 3.550 0.950 3.950 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.450 4.200 1.950 4.600 ;
    END
  END A1
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.200 3.550 2.700 3.950 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.360000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.850 4.850 3.350 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.712500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.900 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.900 8.300 ;
        RECT 0.650 5.550 0.900 7.600 ;
        RECT 2.950 5.550 3.200 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.480000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 0.700 1.600 1.600 ;
        RECT 0.000 0.000 3.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.100 5.200 2.350 7.250 ;
        RECT 2.100 4.900 3.350 5.200 ;
        RECT 1.450 4.250 1.950 4.550 ;
        RECT 0.450 3.600 0.950 3.900 ;
        RECT 2.200 3.600 2.700 3.900 ;
        RECT 2.950 2.600 3.200 4.900 ;
        RECT 2.950 2.350 3.300 2.600 ;
        RECT 0.500 1.850 2.450 2.100 ;
        RECT 0.500 1.050 0.750 1.850 ;
        RECT 2.200 1.050 2.450 1.850 ;
        RECT 3.050 1.050 3.300 2.350 ;
      LAYER Via1 ;
        RECT 2.950 4.900 3.250 5.200 ;
        RECT 1.550 4.250 1.850 4.550 ;
        RECT 0.550 3.600 0.850 3.900 ;
        RECT 2.300 3.600 2.600 3.900 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai21_1


MACRO gf180mcu_osu_sc_gp12t3v3__lshifup
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifup ;
  SIZE 7.800 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 1.020000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 2.600 1.100 2.650 ;
        RECT 4.000 2.600 4.500 2.650 ;
        RECT 0.600 2.300 4.500 2.600 ;
        RECT 0.600 2.250 1.100 2.300 ;
        RECT 4.000 2.250 4.500 2.300 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 6.850 4.200 7.350 4.600 ;
    END
  END Y
  PIN VDDH
    ANTENNADIFFAREA 3.305000 ;
    PORT
      LAYER Nwell ;
        RECT 2.900 5.100 7.800 8.300 ;
      LAYER Metal1 ;
        RECT 2.900 7.600 7.800 8.300 ;
        RECT 4.350 5.550 4.650 7.600 ;
        RECT 6.050 5.550 6.350 7.600 ;
    END
  END VDDH
  PIN VDD
    ANTENNADIFFAREA 1.272500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 2.300 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 2.300 8.300 ;
        RECT 0.550 5.550 0.850 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 3.470000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.850 1.900 ;
        RECT 4.350 0.700 4.650 1.900 ;
        RECT 6.050 0.700 6.350 1.900 ;
        RECT 0.000 0.000 7.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.450 3.300 1.750 7.250 ;
        RECT 3.450 5.200 3.750 7.250 ;
        RECT 4.550 5.200 5.000 5.300 ;
        RECT 3.450 4.900 5.000 5.200 ;
        RECT 1.350 3.000 1.850 3.300 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 1.450 1.050 1.750 3.000 ;
        RECT 3.450 1.050 3.750 4.900 ;
        RECT 4.550 4.850 5.000 4.900 ;
        RECT 5.250 4.550 5.550 7.250 ;
        RECT 6.100 4.900 6.600 5.200 ;
        RECT 6.950 4.550 7.250 7.250 ;
        RECT 4.800 4.100 5.550 4.550 ;
        RECT 6.900 4.250 7.300 4.550 ;
        RECT 4.500 3.000 5.000 3.300 ;
        RECT 4.000 2.300 4.500 2.600 ;
        RECT 5.250 1.050 5.550 4.100 ;
        RECT 6.950 1.050 7.250 4.250 ;
      LAYER Via1 ;
        RECT 4.600 4.900 4.900 5.200 ;
        RECT 1.450 3.000 1.750 3.300 ;
        RECT 0.700 2.300 1.000 2.600 ;
        RECT 6.200 4.900 6.500 5.200 ;
        RECT 6.950 4.250 7.250 4.550 ;
        RECT 4.600 3.000 4.900 3.300 ;
        RECT 4.100 2.300 4.400 2.600 ;
      LAYER Metal2 ;
        RECT 4.550 5.200 4.950 5.250 ;
        RECT 6.100 5.200 6.600 5.250 ;
        RECT 4.500 4.900 6.600 5.200 ;
        RECT 4.550 4.850 4.950 4.900 ;
        RECT 6.100 4.850 6.600 4.900 ;
        RECT 1.350 3.300 1.850 3.350 ;
        RECT 4.500 3.300 5.000 3.350 ;
        RECT 1.350 3.000 5.000 3.300 ;
        RECT 1.350 2.950 1.850 3.000 ;
        RECT 4.500 2.950 5.000 3.000 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifup


MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_4 ;
  SIZE 4.800 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 3.550 0.900 3.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.805000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.950 4.450 3.450 4.850 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.647500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 4.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 4.800 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
        RECT 3.950 5.550 4.200 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.330000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 0.000 0.000 4.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.800 1.650 7.250 ;
        RECT 3.100 4.800 3.350 7.250 ;
        RECT 1.400 4.550 3.350 4.800 ;
        RECT 0.400 3.600 0.900 3.900 ;
        RECT 1.400 2.400 1.650 4.550 ;
        RECT 2.950 4.450 3.350 4.550 ;
        RECT 3.100 2.400 3.350 4.450 ;
        RECT 1.400 2.150 3.350 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
      LAYER Via1 ;
        RECT 0.500 3.600 0.800 3.900 ;
        RECT 3.050 4.500 3.350 4.800 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkinv_4


MACRO gf180mcu_osu_sc_gp12t3v3__inv_4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_4 ;
  SIZE 4.800 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 3.550 0.900 3.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.805000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.950 4.200 3.450 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.647500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 4.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 4.800 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
        RECT 3.950 5.550 4.200 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.330000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 0.000 0.000 4.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.800 1.650 7.250 ;
        RECT 3.100 4.800 3.350 7.250 ;
        RECT 1.400 4.550 3.350 4.800 ;
        RECT 0.400 3.600 0.900 3.900 ;
        RECT 1.400 2.400 1.650 4.550 ;
        RECT 2.950 4.200 3.350 4.550 ;
        RECT 3.100 2.400 3.350 4.200 ;
        RECT 1.400 2.150 3.350 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
      LAYER Via1 ;
        RECT 0.500 3.600 0.800 3.900 ;
        RECT 3.050 4.250 3.350 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__inv_4


MACRO gf180mcu_osu_sc_gp12t3v3__nor2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nor2_1 ;
  SIZE 2.800 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.450 3.550 0.950 3.950 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.850 2.900 2.350 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.317500 ;
    PORT
      LAYER Metal2 ;
        RECT 1.150 4.200 1.650 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 2.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 2.800 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 0.700 0.650 1.900 ;
        RECT 2.100 0.700 2.350 1.900 ;
        RECT 0.000 0.000 2.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.950 5.100 2.200 7.250 ;
        RECT 1.250 4.850 2.200 5.100 ;
        RECT 1.250 4.550 1.500 4.850 ;
        RECT 1.150 4.250 1.650 4.550 ;
        RECT 0.450 3.600 0.950 3.900 ;
        RECT 1.250 1.050 1.500 4.250 ;
        RECT 1.850 2.950 2.350 3.250 ;
      LAYER Via1 ;
        RECT 1.250 4.250 1.550 4.550 ;
        RECT 0.550 3.600 0.850 3.900 ;
        RECT 1.950 2.950 2.250 3.250 ;
  END
END gf180mcu_osu_sc_gp12t3v3__nor2_1


MACRO gf180mcu_osu_sc_gp12t3v3__inv_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_8 ;
  SIZE 8.150 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 6.120000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 3.550 0.900 3.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 5.610001 ;
    PORT
      LAYER Metal2 ;
        RECT 6.350 4.200 6.850 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 6.530001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 8.150 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 8.150 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
        RECT 3.950 5.550 4.200 7.600 ;
        RECT 5.650 5.550 5.900 7.600 ;
        RECT 7.350 5.550 7.600 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.277500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 5.650 0.700 5.900 1.900 ;
        RECT 7.350 0.700 7.600 1.900 ;
        RECT 0.000 0.000 8.150 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.800 1.650 7.250 ;
        RECT 3.100 4.800 3.350 7.250 ;
        RECT 4.800 4.800 5.050 7.250 ;
        RECT 6.500 4.800 6.750 7.250 ;
        RECT 1.400 4.550 6.750 4.800 ;
        RECT 0.400 3.600 0.900 3.900 ;
        RECT 1.400 2.400 1.650 4.550 ;
        RECT 3.100 2.400 3.350 4.550 ;
        RECT 4.800 2.400 5.050 4.550 ;
        RECT 6.350 4.200 6.750 4.550 ;
        RECT 6.500 2.400 6.750 4.200 ;
        RECT 1.400 2.150 6.750 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
        RECT 4.800 1.050 5.050 2.150 ;
        RECT 6.500 1.050 6.750 2.150 ;
      LAYER Via1 ;
        RECT 0.500 3.600 0.800 3.900 ;
        RECT 6.450 4.250 6.750 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__inv_8


MACRO gf180mcu_osu_sc_gp12t3v3__fill_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_16 ;
  SIZE 1.600 BY 8.300 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.600 1.600 8.300 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 1.600 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 5.100 1.600 8.300 ;
  END
END gf180mcu_osu_sc_gp12t3v3__fill_16


MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_2 ;
  SIZE 3.900 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 4.550 1.500 4.600 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 1.100 4.200 1.500 4.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 2.150 4.900 2.650 5.300 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.460000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.900 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.900 8.300 ;
        RECT 1.400 5.550 1.650 7.600 ;
        RECT 3.100 5.550 3.350 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.567500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 0.000 0.000 3.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.300 0.800 7.250 ;
        RECT 2.250 5.250 2.500 7.250 ;
        RECT 2.150 4.950 2.650 5.250 ;
        RECT 1.050 4.250 1.550 4.550 ;
        RECT 0.550 3.000 2.000 3.300 ;
        RECT 0.550 1.050 0.800 3.000 ;
        RECT 2.250 1.050 2.500 4.950 ;
      LAYER Via1 ;
        RECT 2.250 4.950 2.550 5.250 ;
        RECT 1.150 4.250 1.450 4.550 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_2


MACRO gf180mcu_osu_sc_gp12t3v3__or2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__or2_1 ;
  SIZE 3.800 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.900 3.550 1.400 3.950 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.650 2.900 2.150 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.950 4.850 3.450 5.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.202500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.800 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.800 8.300 ;
        RECT 1.950 5.550 2.350 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.905000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 0.700 0.650 1.900 ;
        RECT 2.100 0.700 2.350 1.900 ;
        RECT 0.000 0.000 3.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 5.600 0.800 7.250 ;
        RECT 0.400 5.350 0.800 5.600 ;
        RECT 0.400 4.550 0.650 5.350 ;
        RECT 2.950 5.200 3.200 7.250 ;
        RECT 2.950 4.900 3.450 5.200 ;
        RECT 0.400 4.250 2.700 4.550 ;
        RECT 0.400 2.550 0.650 4.250 ;
        RECT 0.900 3.600 1.400 3.900 ;
        RECT 1.650 2.950 2.150 3.250 ;
        RECT 0.400 2.300 1.500 2.550 ;
        RECT 1.250 1.050 1.500 2.300 ;
        RECT 2.950 1.050 3.200 4.900 ;
      LAYER Via1 ;
        RECT 3.050 4.900 3.350 5.200 ;
        RECT 2.300 4.250 2.600 4.550 ;
        RECT 1.000 3.600 1.300 3.900 ;
        RECT 1.750 2.950 2.050 3.250 ;
      LAYER Metal2 ;
        RECT 2.200 4.200 2.700 4.600 ;
  END
END gf180mcu_osu_sc_gp12t3v3__or2_1


MACRO gf180mcu_osu_sc_gp12t3v3__and2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__and2_1 ;
  SIZE 3.900 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 3.550 1.100 3.950 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.900 2.900 2.400 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.100 4.900 3.600 5.300 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.797500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 3.900 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 3.900 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.607500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.700 2.500 1.900 ;
        RECT 0.000 0.000 3.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.550 1.650 7.250 ;
        RECT 3.100 5.300 3.350 7.250 ;
        RECT 3.100 5.250 3.450 5.300 ;
        RECT 3.100 4.950 3.600 5.250 ;
        RECT 3.100 4.900 3.500 4.950 ;
        RECT 1.300 4.250 2.850 4.550 ;
        RECT 0.600 3.600 1.100 3.900 ;
        RECT 1.400 2.250 1.650 4.250 ;
        RECT 1.900 2.950 2.400 3.250 ;
        RECT 0.700 2.000 1.650 2.250 ;
        RECT 0.700 1.050 0.950 2.000 ;
        RECT 3.100 1.050 3.350 4.900 ;
      LAYER Via1 ;
        RECT 3.200 4.950 3.500 5.250 ;
        RECT 1.400 4.250 1.700 4.550 ;
        RECT 2.450 4.250 2.750 4.550 ;
        RECT 0.700 3.600 1.000 3.900 ;
        RECT 2.000 2.950 2.300 3.250 ;
      LAYER Metal2 ;
        RECT 1.300 4.200 1.800 4.600 ;
        RECT 2.350 4.200 2.850 4.600 ;
  END
END gf180mcu_osu_sc_gp12t3v3__and2_1


MACRO gf180mcu_osu_sc_gp12t3v3__tiel
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tiel ;
  SIZE 2.200 BY 8.300 ;
  PIN Y
    ANTENNADIFFAREA 0.425000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 2.150 1.800 2.550 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 2.200 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 2.200 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.762500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 5.200 1.650 7.250 ;
        RECT 1.150 4.950 1.650 5.200 ;
        RECT 1.400 2.500 1.650 2.550 ;
        RECT 1.300 2.200 1.800 2.500 ;
        RECT 1.400 1.050 1.650 2.200 ;
      LAYER Via1 ;
        RECT 1.400 2.200 1.700 2.500 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tiel


MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_16 ;
  SIZE 15.000 BY 8.300 ;
  PIN A
    ANTENNAGATEAREA 12.240001 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 3.550 0.900 3.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 11.220001 ;
    PORT
      LAYER Metal2 ;
        RECT 13.150 4.450 13.650 4.850 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 12.295001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 5.100 15.000 8.300 ;
      LAYER Metal1 ;
        RECT 0.000 7.600 15.000 8.300 ;
        RECT 0.550 5.550 0.800 7.600 ;
        RECT 2.250 5.550 2.500 7.600 ;
        RECT 3.950 5.550 4.200 7.600 ;
        RECT 5.650 5.550 5.900 7.600 ;
        RECT 7.350 5.550 7.600 7.600 ;
        RECT 9.050 5.550 9.300 7.600 ;
        RECT 10.750 5.550 11.000 7.600 ;
        RECT 12.450 5.550 12.700 7.600 ;
        RECT 14.150 5.550 14.400 7.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.172501 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 5.650 0.700 5.900 1.900 ;
        RECT 7.350 0.700 7.600 1.900 ;
        RECT 9.050 0.700 9.300 1.900 ;
        RECT 10.750 0.700 11.000 1.900 ;
        RECT 12.450 0.700 12.700 1.900 ;
        RECT 14.150 0.700 14.400 1.900 ;
        RECT 0.000 0.000 15.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 4.800 1.650 7.250 ;
        RECT 3.100 4.800 3.350 7.250 ;
        RECT 4.800 4.800 5.050 7.250 ;
        RECT 6.500 4.800 6.750 7.250 ;
        RECT 8.200 4.800 8.450 7.250 ;
        RECT 9.900 4.800 10.150 7.250 ;
        RECT 11.600 4.800 11.850 7.250 ;
        RECT 13.300 4.800 13.550 7.250 ;
        RECT 1.400 4.550 13.550 4.800 ;
        RECT 0.400 3.600 0.900 3.900 ;
        RECT 1.400 2.400 1.650 4.550 ;
        RECT 3.100 2.400 3.350 4.550 ;
        RECT 4.800 2.400 5.050 4.550 ;
        RECT 6.500 2.400 6.750 4.550 ;
        RECT 8.200 2.400 8.450 4.550 ;
        RECT 9.900 2.400 10.150 4.550 ;
        RECT 11.600 2.400 11.850 4.550 ;
        RECT 13.150 4.450 13.550 4.550 ;
        RECT 13.300 2.400 13.550 4.450 ;
        RECT 1.400 2.150 13.550 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
        RECT 4.800 1.050 5.050 2.150 ;
        RECT 6.500 1.050 6.750 2.150 ;
        RECT 8.200 1.050 8.450 2.150 ;
        RECT 9.900 1.050 10.150 2.150 ;
        RECT 11.600 1.050 11.850 2.150 ;
        RECT 13.300 1.050 13.550 2.150 ;
      LAYER Via1 ;
        RECT 0.500 3.600 0.800 3.900 ;
        RECT 13.250 4.500 13.550 4.800 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkinv_16


MACRO gf180mcu_osu_sc_gp12t3v3__fill_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_2 ;
  SIZE 0.900 BY 8.200 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.600 0.200 8.200 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 0.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 5.100 0.200 8.200 ;
  END
END gf180mcu_osu_sc_gp12t3v3__fill_2


END LIBRARY