VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__fill_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_8 ;
  SIZE 0.900 BY 6.350 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.650 0.800 6.350 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 0.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 3.150 0.800 6.350 ;
  END
END gf180mcu_osu_sc_gp9t3v3__fill_8


MACRO gf180mcu_osu_sc_gp9t3v3__oai31_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai31_1 ;
  SIZE 4.900 BY 6.350 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.750 2.250 2.250 2.650 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.550 2.900 3.050 3.300 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.750 2.250 1.250 2.650 ;
    END
  END A2
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.250 2.250 3.750 2.650 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.950 3.900 4.350 3.950 ;
        RECT 3.900 3.600 4.400 3.900 ;
        RECT 3.950 3.550 4.350 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.067500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 4.900 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 4.900 6.350 ;
        RECT 1.000 3.600 1.250 5.650 ;
        RECT 3.950 4.550 4.200 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.242500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.500 ;
        RECT 0.000 0.000 4.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.000 3.900 3.350 5.300 ;
        RECT 3.000 3.600 4.400 3.900 ;
        RECT 4.000 3.550 4.350 3.600 ;
        RECT 2.550 2.950 3.050 3.250 ;
        RECT 0.750 2.300 1.250 2.600 ;
        RECT 1.750 2.300 2.250 2.600 ;
        RECT 3.250 2.300 3.750 2.600 ;
        RECT 1.400 1.750 3.450 2.000 ;
        RECT 1.400 1.050 1.650 1.750 ;
        RECT 3.100 1.050 3.450 1.750 ;
        RECT 4.050 1.050 4.300 3.550 ;
      LAYER Via1 ;
        RECT 4.000 3.600 4.300 3.900 ;
        RECT 2.650 2.950 2.950 3.250 ;
        RECT 0.850 2.300 1.150 2.600 ;
        RECT 1.850 2.300 2.150 2.600 ;
        RECT 3.350 2.300 3.650 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai31_1


MACRO gf180mcu_osu_sc_gp9t3v3__decap_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__decap_1 ;
  SIZE 2.200 BY 6.350 ;
  PIN VDD
    ANTENNADIFFAREA 2.037500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 2.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 2.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 1.400 3.600 1.650 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
END gf180mcu_osu_sc_gp9t3v3__decap_1


MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_2 ;
  SIZE 3.900 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 2.600 1.500 2.650 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 1.100 2.250 1.500 2.300 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 2.150 3.550 2.650 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.797500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.900 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.900 6.350 ;
        RECT 1.400 3.600 1.650 5.650 ;
        RECT 3.100 3.600 3.350 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.905000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 0.000 0.000 3.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.350 0.800 5.300 ;
        RECT 2.250 3.900 2.500 5.300 ;
        RECT 2.150 3.600 2.650 3.900 ;
        RECT 0.550 3.050 2.000 3.350 ;
        RECT 0.550 1.050 0.800 3.050 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 2.250 1.050 2.500 3.600 ;
      LAYER Via1 ;
        RECT 2.250 3.600 2.550 3.900 ;
        RECT 1.150 2.300 1.450 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_2


MACRO gf180mcu_osu_sc_gp9t3v3__tieh
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tieh ;
  SIZE 2.200 BY 6.350 ;
  PIN Y
    ANTENNADIFFAREA 0.850000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 3.550 1.800 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 2.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 2.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.762500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.900 1.650 5.300 ;
        RECT 1.300 3.600 1.800 3.900 ;
        RECT 1.400 3.550 1.650 3.600 ;
        RECT 1.150 2.300 1.650 2.550 ;
        RECT 1.400 1.050 1.650 2.300 ;
      LAYER Via1 ;
        RECT 1.400 3.600 1.700 3.900 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tieh


MACRO gf180mcu_osu_sc_gp9t3v3__xnor2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__xnor2_1 ;
  SIZE 6.400 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.600 3.450 3.950 3.500 ;
        RECT 3.550 3.050 4.000 3.450 ;
        RECT 3.600 3.000 4.000 3.050 ;
        RECT 1.350 2.650 1.650 2.700 ;
        RECT 1.300 2.250 1.700 2.650 ;
        RECT 1.350 1.300 1.650 2.250 ;
        RECT 3.700 1.300 4.000 3.000 ;
        RECT 1.350 1.000 4.000 1.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 4.650 2.650 4.950 2.700 ;
        RECT 4.600 2.600 5.000 2.650 ;
        RECT 4.550 2.300 5.050 2.600 ;
        RECT 4.600 2.250 5.000 2.300 ;
        RECT 4.650 2.200 4.950 2.250 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 2.192500 ;
    PORT
      LAYER Metal2 ;
        RECT 3.000 4.600 3.300 4.850 ;
        RECT 2.950 4.200 3.350 4.600 ;
        RECT 2.950 4.150 3.300 4.200 ;
        RECT 2.950 2.000 3.250 4.150 ;
        RECT 2.900 1.600 3.400 2.000 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.557500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 6.400 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 6.400 6.350 ;
        RECT 1.400 4.700 1.650 5.650 ;
        RECT 4.700 4.700 4.950 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.622500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 4.700 0.700 4.950 1.900 ;
        RECT 0.000 0.000 6.400 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.400 0.800 5.300 ;
        RECT 3.050 4.850 3.300 5.300 ;
        RECT 3.000 4.150 3.300 4.850 ;
        RECT 5.550 3.900 5.800 5.300 ;
        RECT 2.750 3.650 5.800 3.900 ;
        RECT 0.550 3.100 2.400 3.400 ;
        RECT 0.550 1.050 0.800 3.100 ;
        RECT 2.100 2.600 2.400 3.100 ;
        RECT 2.750 3.000 3.050 3.650 ;
        RECT 3.500 3.100 4.000 3.400 ;
        RECT 1.250 2.300 1.750 2.600 ;
        RECT 2.100 2.300 3.500 2.600 ;
        RECT 4.550 2.300 5.050 2.600 ;
        RECT 3.000 1.500 3.300 2.050 ;
        RECT 3.050 1.050 3.300 1.500 ;
        RECT 5.550 1.050 5.800 3.650 ;
      LAYER Via1 ;
        RECT 3.000 4.250 3.300 4.550 ;
        RECT 3.600 3.100 3.900 3.400 ;
        RECT 1.350 2.300 1.650 2.600 ;
        RECT 4.650 2.300 4.950 2.600 ;
        RECT 3.000 1.650 3.300 1.950 ;
  END
END gf180mcu_osu_sc_gp9t3v3__xnor2_1


MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_4 ;
  SIZE 4.800 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 2.250 0.900 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.805000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.300 3.900 3.700 3.950 ;
        RECT 3.250 3.600 3.750 3.900 ;
        RECT 3.300 3.550 3.700 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.732500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 4.800 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 4.800 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.250 3.600 2.500 5.650 ;
        RECT 4.000 3.600 4.250 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.330000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 0.000 0.000 4.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.350 1.650 5.300 ;
        RECT 3.100 3.900 3.350 5.300 ;
        RECT 3.100 3.600 3.750 3.900 ;
        RECT 3.100 3.350 3.350 3.600 ;
        RECT 1.400 3.100 3.350 3.350 ;
        RECT 0.400 2.300 0.900 2.600 ;
        RECT 1.400 2.400 1.650 3.100 ;
        RECT 3.100 2.400 3.350 3.100 ;
        RECT 1.400 2.150 3.350 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
      LAYER Via1 ;
        RECT 3.350 3.600 3.650 3.900 ;
        RECT 0.500 2.300 0.800 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkinv_4


MACRO gf180mcu_osu_sc_gp9t3v3__or2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__or2_1 ;
  SIZE 3.800 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.900 2.250 1.400 2.650 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.650 2.900 2.150 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.950 3.550 3.450 3.950 ;
        RECT 3.050 1.900 3.350 3.550 ;
        RECT 2.950 1.500 3.450 1.900 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.202500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.800 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.800 6.350 ;
        RECT 1.950 4.400 2.350 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.905000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 0.700 0.650 1.550 ;
        RECT 2.100 0.700 2.350 1.900 ;
        RECT 0.000 0.000 3.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.150 0.800 5.300 ;
        RECT 0.550 3.850 2.700 4.150 ;
        RECT 0.550 3.350 0.800 3.850 ;
        RECT 0.400 3.050 0.800 3.350 ;
        RECT 2.400 3.350 2.700 3.850 ;
        RECT 2.950 3.900 3.200 5.300 ;
        RECT 2.950 3.600 3.450 3.900 ;
        RECT 0.400 2.050 0.650 3.050 ;
        RECT 1.650 2.950 2.150 3.250 ;
        RECT 2.400 3.050 2.950 3.350 ;
        RECT 0.900 2.300 1.400 2.600 ;
        RECT 0.400 1.800 1.500 2.050 ;
        RECT 1.250 1.050 1.500 1.800 ;
        RECT 2.950 1.850 3.200 1.900 ;
        RECT 2.950 1.550 3.450 1.850 ;
        RECT 2.950 1.050 3.200 1.550 ;
      LAYER Via1 ;
        RECT 3.050 3.600 3.350 3.900 ;
        RECT 1.750 2.950 2.050 3.250 ;
        RECT 1.000 2.300 1.300 2.600 ;
        RECT 3.050 1.550 3.350 1.850 ;
  END
END gf180mcu_osu_sc_gp9t3v3__or2_1


MACRO gf180mcu_osu_sc_gp9t3v3__inv_4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_4 ;
  SIZE 4.800 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 2.250 0.900 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.805000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.300 3.900 3.700 3.950 ;
        RECT 3.250 3.600 3.750 3.900 ;
        RECT 3.300 3.550 3.700 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.732500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 4.800 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 4.800 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.250 3.600 2.500 5.650 ;
        RECT 4.000 3.600 4.250 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.330000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 0.000 0.000 4.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.350 1.650 5.300 ;
        RECT 3.100 3.900 3.350 5.300 ;
        RECT 3.100 3.600 3.750 3.900 ;
        RECT 3.100 3.350 3.350 3.600 ;
        RECT 1.400 3.100 3.350 3.350 ;
        RECT 0.400 2.300 0.900 2.600 ;
        RECT 1.400 2.400 1.650 3.100 ;
        RECT 3.100 2.400 3.350 3.100 ;
        RECT 1.400 2.150 3.350 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
      LAYER Via1 ;
        RECT 3.350 3.600 3.650 3.900 ;
        RECT 0.500 2.300 0.800 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__inv_4


MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_1 ;
  SIZE 2.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.550 2.250 1.050 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 3.550 1.800 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 2.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 2.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.762500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.900 1.650 5.300 ;
        RECT 1.300 3.600 1.800 3.900 ;
        RECT 0.550 2.300 1.050 2.600 ;
        RECT 1.400 1.050 1.650 3.600 ;
      LAYER Via1 ;
        RECT 1.400 3.600 1.700 3.900 ;
        RECT 0.650 2.300 0.950 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkinv_1


MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_8 ;
  SIZE 9.050 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 2.600 1.500 2.650 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 1.100 2.250 1.500 2.300 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 5.610001 ;
    PORT
      LAYER Metal2 ;
        RECT 7.250 3.550 7.750 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 6.952500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 9.050 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 9.050 6.350 ;
        RECT 1.400 3.600 1.650 5.650 ;
        RECT 3.100 3.600 3.350 5.650 ;
        RECT 4.800 3.600 5.050 5.650 ;
        RECT 6.500 3.600 6.750 5.650 ;
        RECT 8.200 3.600 8.450 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.657500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.900 ;
        RECT 8.200 0.700 8.450 1.900 ;
        RECT 0.000 0.000 9.050 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.350 0.800 5.300 ;
        RECT 2.250 3.350 2.500 5.300 ;
        RECT 3.950 3.350 4.200 5.300 ;
        RECT 5.650 3.350 5.900 5.300 ;
        RECT 7.350 3.900 7.600 5.300 ;
        RECT 7.250 3.600 7.750 3.900 ;
        RECT 7.350 3.350 7.600 3.600 ;
        RECT 0.550 3.050 2.000 3.350 ;
        RECT 2.250 3.050 7.600 3.350 ;
        RECT 0.550 1.050 0.800 3.050 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 2.250 2.450 2.500 3.050 ;
        RECT 3.950 2.450 4.200 3.050 ;
        RECT 5.650 2.450 5.900 3.050 ;
        RECT 7.350 2.450 7.600 3.050 ;
        RECT 2.250 2.150 7.600 2.450 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
        RECT 5.650 1.050 5.900 2.150 ;
        RECT 7.350 1.050 7.600 2.150 ;
      LAYER Via1 ;
        RECT 7.350 3.600 7.650 3.900 ;
        RECT 1.150 2.300 1.450 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_8


MACRO gf180mcu_osu_sc_gp9t3v3__inv_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_8 ;
  SIZE 8.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 6.120000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 2.250 0.900 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 5.610001 ;
    PORT
      LAYER Metal2 ;
        RECT 6.700 3.900 7.100 3.950 ;
        RECT 6.650 3.600 7.150 3.900 ;
        RECT 6.700 3.550 7.100 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 6.615000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 8.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 8.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.250 3.600 2.500 5.650 ;
        RECT 3.950 3.600 4.200 5.650 ;
        RECT 5.650 3.600 5.900 5.650 ;
        RECT 7.400 3.600 7.650 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.277500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 5.650 0.700 5.900 1.900 ;
        RECT 7.350 0.700 7.600 1.900 ;
        RECT 0.000 0.000 8.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.350 1.650 5.300 ;
        RECT 3.100 3.350 3.350 5.300 ;
        RECT 4.800 3.350 5.050 5.300 ;
        RECT 6.500 3.900 6.750 5.300 ;
        RECT 6.500 3.600 7.150 3.900 ;
        RECT 6.500 3.350 6.750 3.600 ;
        RECT 1.400 3.100 6.750 3.350 ;
        RECT 0.400 2.300 0.900 2.600 ;
        RECT 1.400 2.400 1.650 3.100 ;
        RECT 3.100 2.400 3.350 3.100 ;
        RECT 4.800 2.400 5.050 3.100 ;
        RECT 6.500 2.400 6.750 3.100 ;
        RECT 1.400 2.150 6.750 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
        RECT 4.800 1.050 5.050 2.150 ;
        RECT 6.500 1.050 6.750 2.150 ;
      LAYER Via1 ;
        RECT 6.750 3.600 7.050 3.900 ;
        RECT 0.500 2.300 0.800 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__inv_8


MACRO gf180mcu_osu_sc_gp9t3v3__mux2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__mux2_1 ;
  SIZE 5.100 BY 6.350 ;
  PIN A
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.350 2.250 2.850 2.650 ;
    END
  END A
  PIN B
    ANTENNADIFFAREA 1.657500 ;
    PORT
      LAYER Metal2 ;
        RECT 4.250 2.250 4.750 2.650 ;
    END
  END B
  PIN Sel
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.550 2.900 1.050 3.300 ;
    END
  END Sel
  PIN Y
    ANTENNADIFFAREA 1.785000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.000 4.200 3.500 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.200000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 5.100 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 5.100 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.775000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 5.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.450 1.650 5.300 ;
        RECT 0.550 2.950 1.050 3.250 ;
        RECT 1.400 3.150 1.950 3.450 ;
        RECT 1.400 2.400 1.650 3.150 ;
        RECT 2.250 2.650 2.500 5.300 ;
        RECT 3.100 4.650 3.350 5.300 ;
        RECT 3.100 4.150 3.400 4.650 ;
        RECT 1.400 2.100 2.000 2.400 ;
        RECT 2.250 2.250 2.850 2.650 ;
        RECT 1.400 1.050 1.650 2.100 ;
        RECT 2.250 1.050 2.500 2.250 ;
        RECT 3.100 1.050 3.350 4.150 ;
        RECT 3.650 3.000 3.950 3.550 ;
        RECT 4.250 2.650 4.500 5.300 ;
        RECT 4.250 2.250 4.750 2.650 ;
        RECT 4.250 1.050 4.500 2.250 ;
      LAYER Via1 ;
        RECT 0.650 2.950 0.950 3.250 ;
        RECT 1.550 3.150 1.850 3.450 ;
        RECT 3.100 4.250 3.400 4.550 ;
        RECT 2.450 2.300 2.750 2.600 ;
        RECT 3.650 3.150 3.950 3.450 ;
        RECT 4.350 2.300 4.650 2.600 ;
      LAYER Metal2 ;
        RECT 1.450 3.450 1.950 3.500 ;
        RECT 3.550 3.450 4.050 3.500 ;
        RECT 1.450 3.150 4.050 3.450 ;
        RECT 1.450 3.100 1.950 3.150 ;
        RECT 3.550 3.100 4.050 3.150 ;
  END
END gf180mcu_osu_sc_gp9t3v3__mux2_1


MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_16 ;
  SIZE 15.800 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 2.600 1.500 2.650 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 1.100 2.250 1.500 2.300 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 11.220001 ;
    PORT
      LAYER Metal2 ;
        RECT 14.050 3.550 14.550 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 12.380001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 15.800 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 15.800 6.350 ;
        RECT 1.400 3.600 1.650 5.650 ;
        RECT 3.100 3.600 3.350 5.650 ;
        RECT 4.800 3.600 5.050 5.650 ;
        RECT 6.500 3.600 6.750 5.650 ;
        RECT 8.200 3.600 8.450 5.650 ;
        RECT 9.900 3.600 10.150 5.650 ;
        RECT 11.600 3.600 11.850 5.650 ;
        RECT 13.300 3.600 13.550 5.650 ;
        RECT 15.000 3.600 15.250 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.215000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.900 ;
        RECT 8.200 0.700 8.450 1.900 ;
        RECT 9.900 0.700 10.150 1.900 ;
        RECT 11.600 0.700 11.850 1.900 ;
        RECT 13.300 0.700 13.550 1.900 ;
        RECT 15.000 0.700 15.250 1.900 ;
        RECT 0.000 0.000 15.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.350 0.800 5.300 ;
        RECT 2.250 3.350 2.500 5.300 ;
        RECT 3.950 3.350 4.200 5.300 ;
        RECT 5.650 3.350 5.900 5.300 ;
        RECT 7.350 3.350 7.600 5.300 ;
        RECT 9.050 3.350 9.300 5.300 ;
        RECT 10.750 3.350 11.000 5.300 ;
        RECT 12.450 3.350 12.700 5.300 ;
        RECT 14.150 3.900 14.400 5.300 ;
        RECT 14.050 3.600 14.550 3.900 ;
        RECT 14.150 3.350 14.400 3.600 ;
        RECT 0.550 3.050 2.000 3.350 ;
        RECT 2.250 3.050 14.400 3.350 ;
        RECT 0.550 1.050 0.800 3.050 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 2.250 2.450 2.500 3.050 ;
        RECT 3.950 2.450 4.200 3.050 ;
        RECT 5.650 2.450 5.900 3.050 ;
        RECT 7.350 2.450 7.600 3.050 ;
        RECT 9.050 2.450 9.300 3.050 ;
        RECT 10.750 2.450 11.000 3.050 ;
        RECT 12.450 2.450 12.700 3.050 ;
        RECT 14.150 2.450 14.400 3.050 ;
        RECT 2.250 2.150 14.400 2.450 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
        RECT 5.650 1.050 5.900 2.150 ;
        RECT 7.350 1.050 7.600 2.150 ;
        RECT 9.050 1.050 9.300 2.150 ;
        RECT 10.750 1.050 11.000 2.150 ;
        RECT 12.450 1.050 12.700 2.150 ;
        RECT 14.150 1.050 14.400 2.150 ;
      LAYER Via1 ;
        RECT 14.150 3.600 14.450 3.900 ;
        RECT 1.150 2.300 1.450 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_16


MACRO gf180mcu_osu_sc_gp9t3v3__dffn_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dffn_1 ;
  SIZE 15.500 BY 6.350 ;
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.750 3.250 2.250 3.300 ;
        RECT 1.700 2.950 2.300 3.250 ;
        RECT 1.750 2.900 2.250 2.950 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.100 3.250 11.500 3.300 ;
        RECT 11.050 2.950 11.550 3.250 ;
        RECT 11.100 2.900 11.500 2.950 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.800 4.550 15.200 4.600 ;
        RECT 14.750 4.250 15.250 4.550 ;
        RECT 14.800 4.200 15.200 4.250 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 0.765000 ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.000 3.900 14.400 3.950 ;
        RECT 13.950 3.600 14.450 3.900 ;
        RECT 14.000 3.550 14.400 3.600 ;
    END
  END QN
  PIN VDD
    ANTENNADIFFAREA 8.725000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 15.500 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 15.500 6.350 ;
        RECT 1.400 4.850 1.650 5.650 ;
        RECT 5.000 4.200 5.250 5.650 ;
        RECT 8.600 4.850 8.850 5.650 ;
        RECT 11.400 3.600 11.650 5.650 ;
        RECT 13.850 4.150 14.100 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 6.312500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.600 ;
        RECT 5.000 0.700 5.250 1.500 ;
        RECT 8.600 0.700 8.850 1.600 ;
        RECT 11.400 0.700 11.650 1.500 ;
        RECT 13.850 0.700 14.100 1.700 ;
        RECT 0.000 0.000 15.500 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.450 0.800 5.300 ;
        RECT 3.300 4.600 3.850 5.300 ;
        RECT 0.500 2.400 0.800 2.450 ;
        RECT 0.400 2.100 0.800 2.400 ;
        RECT 0.500 2.000 0.800 2.100 ;
        RECT 0.550 1.050 0.800 2.000 ;
        RECT 1.050 4.300 3.850 4.600 ;
        RECT 1.050 3.400 1.350 4.300 ;
        RECT 6.400 4.200 6.950 5.300 ;
        RECT 8.050 4.300 8.550 4.600 ;
        RECT 8.150 4.200 8.450 4.300 ;
        RECT 9.450 4.100 9.700 5.300 ;
        RECT 2.650 3.650 8.900 3.950 ;
        RECT 9.450 3.850 10.000 4.100 ;
        RECT 2.650 3.400 2.950 3.650 ;
        RECT 1.050 3.100 1.450 3.400 ;
        RECT 1.050 2.150 1.350 3.100 ;
        RECT 1.750 2.950 2.250 3.250 ;
        RECT 2.500 3.100 2.950 3.400 ;
        RECT 2.650 3.050 2.950 3.100 ;
        RECT 4.700 2.400 5.000 2.450 ;
        RECT 1.050 1.900 2.250 2.150 ;
        RECT 2.700 2.100 3.200 2.400 ;
        RECT 4.600 2.100 5.100 2.400 ;
        RECT 6.050 2.350 6.350 3.650 ;
        RECT 8.600 3.400 8.900 3.650 ;
        RECT 8.600 3.250 9.450 3.400 ;
        RECT 8.600 3.100 9.500 3.250 ;
        RECT 7.250 3.000 7.550 3.050 ;
        RECT 7.200 2.600 7.600 3.000 ;
        RECT 9.000 2.950 9.500 3.100 ;
        RECT 9.750 2.600 10.000 3.850 ;
        RECT 10.550 3.300 10.800 5.300 ;
        RECT 10.500 3.250 10.800 3.300 ;
        RECT 10.250 2.950 10.800 3.250 ;
        RECT 10.500 2.900 10.800 2.950 ;
        RECT 7.250 2.550 7.550 2.600 ;
        RECT 5.950 2.050 6.450 2.350 ;
        RECT 8.050 2.300 8.550 2.600 ;
        RECT 9.450 2.300 10.000 2.600 ;
        RECT 2.000 1.750 2.250 1.900 ;
        RECT 2.000 1.500 3.850 1.750 ;
        RECT 3.300 1.050 3.850 1.500 ;
        RECT 6.400 1.050 6.950 1.750 ;
        RECT 7.250 1.550 7.550 2.050 ;
        RECT 9.450 1.550 9.750 2.300 ;
        RECT 9.450 1.050 9.700 1.550 ;
        RECT 10.550 1.050 10.800 2.900 ;
        RECT 11.150 2.850 11.450 3.350 ;
        RECT 12.250 2.950 12.500 5.300 ;
        RECT 13.000 3.900 13.250 5.300 ;
        RECT 14.700 4.600 14.950 5.300 ;
        RECT 14.700 4.250 15.250 4.600 ;
        RECT 14.700 4.200 15.200 4.250 ;
        RECT 13.000 3.600 14.450 3.900 ;
        RECT 12.250 2.650 13.650 2.950 ;
        RECT 11.600 2.050 11.900 2.550 ;
        RECT 11.500 1.750 12.000 2.050 ;
        RECT 12.250 1.050 12.500 2.650 ;
        RECT 14.050 2.200 14.350 3.600 ;
        RECT 13.000 1.950 14.350 2.200 ;
        RECT 13.000 1.050 13.250 1.950 ;
        RECT 14.700 1.050 14.950 4.200 ;
      LAYER Via1 ;
        RECT 0.500 2.100 0.800 2.400 ;
        RECT 6.500 4.300 6.800 4.600 ;
        RECT 8.150 4.300 8.450 4.600 ;
        RECT 1.850 2.950 2.150 3.250 ;
        RECT 2.800 2.100 3.100 2.400 ;
        RECT 4.700 2.100 5.000 2.400 ;
        RECT 9.100 2.950 9.400 3.250 ;
        RECT 7.250 2.650 7.550 2.950 ;
        RECT 10.350 2.950 10.650 3.250 ;
        RECT 8.150 2.300 8.450 2.600 ;
        RECT 6.500 1.450 6.800 1.750 ;
        RECT 7.250 1.650 7.550 1.950 ;
        RECT 9.450 1.650 9.750 1.950 ;
        RECT 11.150 2.950 11.450 3.250 ;
        RECT 14.850 4.250 15.150 4.550 ;
        RECT 14.050 3.600 14.350 3.900 ;
        RECT 13.250 2.650 13.550 2.950 ;
        RECT 11.600 1.750 11.900 2.050 ;
      LAYER Metal2 ;
        RECT 2.800 5.000 7.550 5.300 ;
        RECT 2.800 2.450 3.100 5.000 ;
        RECT 6.500 4.650 6.800 4.700 ;
        RECT 6.450 4.250 6.850 4.650 ;
        RECT 0.450 2.400 0.850 2.450 ;
        RECT 2.750 2.400 3.200 2.450 ;
        RECT 4.650 2.400 5.050 2.450 ;
        RECT 0.400 2.100 0.900 2.400 ;
        RECT 2.700 2.100 3.200 2.400 ;
        RECT 4.600 2.100 5.100 2.400 ;
        RECT 0.450 2.050 0.850 2.100 ;
        RECT 2.750 2.050 3.200 2.100 ;
        RECT 4.650 2.050 5.050 2.100 ;
        RECT 0.500 1.450 0.800 2.050 ;
        RECT 4.700 1.450 5.000 2.050 ;
        RECT 6.500 1.800 6.800 4.250 ;
        RECT 7.250 3.800 7.550 5.000 ;
        RECT 8.100 4.600 8.500 4.650 ;
        RECT 8.050 4.300 12.450 4.600 ;
        RECT 8.100 4.250 8.500 4.300 ;
        RECT 7.200 3.500 7.550 3.800 ;
        RECT 7.200 3.050 7.500 3.500 ;
        RECT 7.200 2.550 7.600 3.050 ;
        RECT 8.150 2.650 8.450 4.250 ;
        RECT 9.050 3.250 9.450 3.300 ;
        RECT 10.300 3.250 10.700 3.300 ;
        RECT 9.000 2.950 10.750 3.250 ;
        RECT 12.150 2.950 12.450 4.300 ;
        RECT 13.200 2.950 13.600 3.000 ;
        RECT 9.050 2.900 9.450 2.950 ;
        RECT 10.300 2.900 10.700 2.950 ;
        RECT 12.150 2.650 13.650 2.950 ;
        RECT 8.100 2.600 8.500 2.650 ;
        RECT 13.200 2.600 13.600 2.650 ;
        RECT 7.250 2.000 7.550 2.550 ;
        RECT 8.050 2.300 8.550 2.600 ;
        RECT 8.100 2.250 8.500 2.300 ;
        RECT 11.550 2.050 11.950 2.100 ;
        RECT 7.200 1.950 7.600 2.000 ;
        RECT 9.400 1.950 9.800 2.000 ;
        RECT 0.500 1.150 5.000 1.450 ;
        RECT 6.450 1.400 6.850 1.800 ;
        RECT 7.150 1.650 9.900 1.950 ;
        RECT 11.200 1.750 12.000 2.050 ;
        RECT 11.200 1.700 11.950 1.750 ;
        RECT 7.200 1.600 7.600 1.650 ;
        RECT 9.400 1.600 9.800 1.650 ;
        RECT 6.500 1.300 6.850 1.400 ;
        RECT 11.200 1.300 11.500 1.700 ;
        RECT 6.500 1.000 11.750 1.300 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dffn_1


MACRO gf180mcu_osu_sc_gp9t3v3__fill_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_2 ;
  SIZE 0.900 BY 6.350 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.650 0.200 6.350 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 0.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 3.150 0.200 6.350 ;
  END
END gf180mcu_osu_sc_gp9t3v3__fill_2


MACRO gf180mcu_osu_sc_gp9t3v3__inv_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_16 ;
  SIZE 15.000 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 12.240001 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 2.250 0.900 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 11.220001 ;
    PORT
      LAYER Metal2 ;
        RECT 13.400 3.900 13.800 3.950 ;
        RECT 13.350 3.600 13.850 3.900 ;
        RECT 13.400 3.550 13.800 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 12.380001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 15.000 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 15.000 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.250 3.600 2.500 5.650 ;
        RECT 3.950 3.600 4.200 5.650 ;
        RECT 5.650 3.600 5.900 5.650 ;
        RECT 7.350 3.600 7.600 5.650 ;
        RECT 9.050 3.600 9.300 5.650 ;
        RECT 10.750 3.600 11.000 5.650 ;
        RECT 12.450 3.600 12.700 5.650 ;
        RECT 14.150 3.600 14.400 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.172501 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 5.650 0.700 5.900 1.900 ;
        RECT 7.350 0.700 7.600 1.900 ;
        RECT 9.050 0.700 9.300 1.900 ;
        RECT 10.750 0.700 11.000 1.900 ;
        RECT 12.450 0.700 12.700 1.900 ;
        RECT 14.150 0.700 14.400 1.900 ;
        RECT 0.000 0.000 15.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.350 1.650 5.300 ;
        RECT 3.100 3.350 3.350 5.300 ;
        RECT 4.800 3.350 5.050 5.300 ;
        RECT 6.500 3.350 6.750 5.300 ;
        RECT 8.200 3.350 8.450 5.300 ;
        RECT 9.900 3.350 10.150 5.300 ;
        RECT 11.600 3.350 11.850 5.300 ;
        RECT 13.300 3.900 13.550 5.300 ;
        RECT 13.300 3.600 13.850 3.900 ;
        RECT 13.300 3.350 13.550 3.600 ;
        RECT 1.400 3.100 13.550 3.350 ;
        RECT 0.400 2.300 0.900 2.600 ;
        RECT 1.400 2.400 1.650 3.100 ;
        RECT 3.100 2.400 3.350 3.100 ;
        RECT 4.800 2.400 5.050 3.100 ;
        RECT 6.500 2.400 6.750 3.100 ;
        RECT 8.200 2.400 8.450 3.100 ;
        RECT 9.900 2.400 10.150 3.100 ;
        RECT 11.600 2.400 11.850 3.100 ;
        RECT 13.300 2.400 13.550 3.100 ;
        RECT 1.400 2.150 13.550 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
        RECT 4.800 1.050 5.050 2.150 ;
        RECT 6.500 1.050 6.750 2.150 ;
        RECT 8.200 1.050 8.450 2.150 ;
        RECT 9.900 1.050 10.150 2.150 ;
        RECT 11.600 1.050 11.850 2.150 ;
        RECT 13.300 1.050 13.550 2.150 ;
      LAYER Via1 ;
        RECT 13.450 3.600 13.750 3.900 ;
        RECT 0.500 2.300 0.800 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__inv_16


MACRO gf180mcu_osu_sc_gp9t3v3__dff_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dff_1 ;
  SIZE 14.500 BY 6.350 ;
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.750 3.250 2.250 3.300 ;
        RECT 1.700 2.950 2.300 3.250 ;
        RECT 1.750 2.900 2.250 2.950 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.050 3.250 9.450 3.300 ;
        RECT 9.000 2.950 9.500 3.250 ;
        RECT 9.050 2.900 9.450 2.950 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.800 4.550 14.200 4.600 ;
        RECT 13.750 4.250 14.250 4.550 ;
        RECT 13.800 4.200 14.200 4.250 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 0.765000 ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.000 3.900 13.400 3.950 ;
        RECT 12.950 3.600 13.450 3.900 ;
        RECT 13.000 3.550 13.400 3.600 ;
    END
  END QN
  PIN VDD
    ANTENNADIFFAREA 8.302501 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 14.500 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 14.500 6.350 ;
        RECT 1.400 4.850 1.650 5.650 ;
        RECT 5.000 4.200 5.250 5.650 ;
        RECT 8.600 4.850 8.850 5.650 ;
        RECT 10.400 3.600 10.650 5.650 ;
        RECT 12.850 4.150 13.100 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 5.932500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.600 ;
        RECT 5.000 0.700 5.250 1.500 ;
        RECT 8.600 0.700 8.850 1.600 ;
        RECT 10.400 0.700 10.650 1.500 ;
        RECT 12.850 0.700 13.100 1.700 ;
        RECT 0.000 0.000 14.500 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.450 0.800 5.300 ;
        RECT 3.300 4.600 3.850 5.300 ;
        RECT 0.500 2.400 0.800 2.450 ;
        RECT 0.400 2.100 0.800 2.400 ;
        RECT 0.500 2.000 0.800 2.100 ;
        RECT 0.550 1.050 0.800 2.000 ;
        RECT 1.050 4.300 3.850 4.600 ;
        RECT 1.050 3.400 1.350 4.300 ;
        RECT 6.400 4.200 6.950 5.300 ;
        RECT 8.050 4.300 8.550 4.600 ;
        RECT 8.150 4.200 8.450 4.300 ;
        RECT 2.650 3.650 8.950 3.950 ;
        RECT 2.650 3.400 2.950 3.650 ;
        RECT 1.050 3.100 1.450 3.400 ;
        RECT 1.050 2.150 1.350 3.100 ;
        RECT 1.750 2.950 2.250 3.250 ;
        RECT 2.500 3.100 3.000 3.400 ;
        RECT 4.700 2.400 5.000 2.450 ;
        RECT 1.050 1.900 2.250 2.150 ;
        RECT 2.700 2.100 3.200 2.400 ;
        RECT 4.600 2.100 5.100 2.400 ;
        RECT 6.050 2.350 6.350 3.650 ;
        RECT 8.650 3.350 8.950 3.650 ;
        RECT 9.450 3.850 9.700 5.300 ;
        RECT 9.450 3.600 10.000 3.850 ;
        RECT 8.650 3.250 9.400 3.350 ;
        RECT 7.200 2.950 7.700 3.250 ;
        RECT 8.650 2.950 9.500 3.250 ;
        RECT 9.750 2.600 10.000 3.600 ;
        RECT 5.950 2.050 6.450 2.350 ;
        RECT 8.050 2.300 8.550 2.600 ;
        RECT 9.450 2.300 10.000 2.600 ;
        RECT 2.000 1.750 2.250 1.900 ;
        RECT 2.000 1.500 3.850 1.750 ;
        RECT 3.300 1.050 3.850 1.500 ;
        RECT 6.400 1.050 6.950 1.750 ;
        RECT 7.250 1.550 7.550 2.050 ;
        RECT 9.450 1.550 9.750 2.300 ;
        RECT 10.600 2.050 10.900 3.050 ;
        RECT 11.250 2.950 11.500 5.300 ;
        RECT 12.000 3.900 12.250 5.300 ;
        RECT 13.700 4.600 13.950 5.300 ;
        RECT 13.700 4.250 14.250 4.600 ;
        RECT 13.700 4.200 14.200 4.250 ;
        RECT 12.000 3.600 13.450 3.900 ;
        RECT 11.250 2.650 12.650 2.950 ;
        RECT 10.500 1.750 11.000 2.050 ;
        RECT 9.450 1.050 9.700 1.550 ;
        RECT 11.250 1.050 11.500 2.650 ;
        RECT 13.050 2.200 13.350 3.600 ;
        RECT 12.000 1.950 13.350 2.200 ;
        RECT 12.000 1.050 12.250 1.950 ;
        RECT 13.700 1.050 13.950 4.200 ;
      LAYER Via1 ;
        RECT 0.500 2.100 0.800 2.400 ;
        RECT 6.500 4.300 6.800 4.600 ;
        RECT 8.150 4.300 8.450 4.600 ;
        RECT 1.850 2.950 2.150 3.250 ;
        RECT 2.800 2.100 3.100 2.400 ;
        RECT 4.700 2.100 5.000 2.400 ;
        RECT 7.300 2.950 7.600 3.250 ;
        RECT 9.100 2.950 9.400 3.250 ;
        RECT 8.150 2.300 8.450 2.600 ;
        RECT 6.500 1.450 6.800 1.750 ;
        RECT 7.250 1.650 7.550 1.950 ;
        RECT 13.850 4.250 14.150 4.550 ;
        RECT 13.050 3.600 13.350 3.900 ;
        RECT 12.250 2.650 12.550 2.950 ;
        RECT 9.450 1.650 9.750 1.950 ;
        RECT 10.600 1.750 10.900 2.050 ;
      LAYER Metal2 ;
        RECT 2.800 5.000 7.550 5.300 ;
        RECT 2.800 2.450 3.100 5.000 ;
        RECT 6.500 4.650 6.800 4.700 ;
        RECT 6.450 4.250 6.850 4.650 ;
        RECT 0.450 2.400 0.850 2.450 ;
        RECT 2.750 2.400 3.200 2.450 ;
        RECT 4.650 2.400 5.050 2.450 ;
        RECT 0.400 2.100 0.900 2.400 ;
        RECT 2.700 2.100 3.200 2.400 ;
        RECT 4.600 2.100 5.100 2.400 ;
        RECT 0.450 2.050 0.850 2.100 ;
        RECT 2.750 2.050 3.200 2.100 ;
        RECT 4.650 2.050 5.050 2.100 ;
        RECT 0.500 1.450 0.800 2.050 ;
        RECT 4.700 1.450 5.000 2.050 ;
        RECT 6.500 1.800 6.800 4.250 ;
        RECT 7.250 3.350 7.550 5.000 ;
        RECT 8.100 4.600 8.500 4.650 ;
        RECT 8.050 4.300 11.450 4.600 ;
        RECT 8.100 4.250 8.500 4.300 ;
        RECT 7.250 2.900 7.650 3.350 ;
        RECT 7.250 2.000 7.550 2.900 ;
        RECT 8.150 2.650 8.450 4.250 ;
        RECT 11.150 2.950 11.450 4.300 ;
        RECT 12.200 2.950 12.600 3.000 ;
        RECT 11.150 2.650 12.650 2.950 ;
        RECT 8.100 2.600 8.500 2.650 ;
        RECT 12.200 2.600 12.600 2.650 ;
        RECT 8.050 2.300 8.550 2.600 ;
        RECT 8.100 2.250 8.500 2.300 ;
        RECT 10.550 2.050 10.950 2.100 ;
        RECT 7.200 1.950 7.600 2.000 ;
        RECT 9.400 1.950 9.800 2.000 ;
        RECT 0.500 1.150 5.000 1.450 ;
        RECT 6.450 1.400 6.850 1.800 ;
        RECT 7.150 1.650 9.900 1.950 ;
        RECT 10.200 1.750 11.000 2.050 ;
        RECT 10.200 1.700 10.950 1.750 ;
        RECT 7.200 1.600 7.600 1.650 ;
        RECT 9.400 1.600 9.800 1.650 ;
        RECT 6.500 1.300 6.850 1.400 ;
        RECT 10.200 1.300 10.500 1.700 ;
        RECT 6.500 1.000 10.500 1.300 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dff_1


MACRO gf180mcu_osu_sc_gp9t3v3__aoi21_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__aoi21_1 ;
  SIZE 3.900 BY 6.350 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 2.250 1.100 2.650 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.600 2.900 2.100 3.300 ;
    END
  END A1
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.350 2.250 2.850 2.650 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.317500 ;
    PORT
      LAYER Metal2 ;
        RECT 3.000 3.550 3.500 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.947500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.900 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.900 6.350 ;
        RECT 1.400 4.350 1.650 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.862500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 0.700 0.950 1.900 ;
        RECT 2.950 0.700 3.200 1.500 ;
        RECT 0.000 0.000 3.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.100 0.800 5.300 ;
        RECT 2.250 4.100 2.500 5.300 ;
        RECT 0.550 3.850 2.500 4.100 ;
        RECT 3.100 3.900 3.350 5.300 ;
        RECT 3.000 3.600 3.500 3.900 ;
        RECT 1.600 2.950 2.100 3.250 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 2.350 2.300 2.850 2.600 ;
        RECT 3.100 2.000 3.350 3.600 ;
        RECT 2.100 1.750 3.350 2.000 ;
        RECT 2.100 1.050 2.350 1.750 ;
      LAYER Via1 ;
        RECT 3.100 3.600 3.400 3.900 ;
        RECT 1.700 2.950 2.000 3.250 ;
        RECT 0.700 2.300 1.000 2.600 ;
        RECT 2.450 2.300 2.750 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__aoi21_1


MACRO gf180mcu_osu_sc_gp9t3v3__buf_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_16 ;
  SIZE 15.800 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 2.600 1.500 2.650 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 1.100 2.250 1.500 2.300 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 11.220001 ;
    PORT
      LAYER Metal2 ;
        RECT 14.050 3.550 14.550 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 12.380001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 15.800 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 15.800 6.350 ;
        RECT 1.400 3.600 1.650 5.650 ;
        RECT 3.100 3.600 3.350 5.650 ;
        RECT 4.800 3.600 5.050 5.650 ;
        RECT 6.500 3.600 6.750 5.650 ;
        RECT 8.200 3.600 8.450 5.650 ;
        RECT 9.900 3.600 10.150 5.650 ;
        RECT 11.600 3.600 11.850 5.650 ;
        RECT 13.300 3.600 13.550 5.650 ;
        RECT 15.000 3.600 15.250 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.215000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.900 ;
        RECT 8.200 0.700 8.450 1.900 ;
        RECT 9.900 0.700 10.150 1.900 ;
        RECT 11.600 0.700 11.850 1.900 ;
        RECT 13.300 0.700 13.550 1.900 ;
        RECT 15.000 0.700 15.250 1.900 ;
        RECT 0.000 0.000 15.800 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.350 0.800 5.300 ;
        RECT 2.250 3.350 2.500 5.300 ;
        RECT 3.950 3.350 4.200 5.300 ;
        RECT 5.650 3.350 5.900 5.300 ;
        RECT 7.350 3.350 7.600 5.300 ;
        RECT 9.050 3.350 9.300 5.300 ;
        RECT 10.750 3.350 11.000 5.300 ;
        RECT 12.450 3.350 12.700 5.300 ;
        RECT 14.150 3.900 14.400 5.300 ;
        RECT 14.050 3.600 14.550 3.900 ;
        RECT 14.150 3.350 14.400 3.600 ;
        RECT 0.550 3.050 2.000 3.350 ;
        RECT 2.250 3.050 14.400 3.350 ;
        RECT 0.550 1.050 0.800 3.050 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 2.250 2.450 2.500 3.050 ;
        RECT 3.950 2.450 4.200 3.050 ;
        RECT 5.650 2.450 5.900 3.050 ;
        RECT 7.350 2.450 7.600 3.050 ;
        RECT 9.050 2.450 9.300 3.050 ;
        RECT 10.750 2.450 11.000 3.050 ;
        RECT 12.450 2.450 12.700 3.050 ;
        RECT 14.150 2.450 14.400 3.050 ;
        RECT 2.250 2.150 14.400 2.450 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
        RECT 5.650 1.050 5.900 2.150 ;
        RECT 7.350 1.050 7.600 2.150 ;
        RECT 9.050 1.050 9.300 2.150 ;
        RECT 10.750 1.050 11.000 2.150 ;
        RECT 12.450 1.050 12.700 2.150 ;
        RECT 14.150 1.050 14.400 2.150 ;
      LAYER Via1 ;
        RECT 14.150 3.600 14.450 3.900 ;
        RECT 1.150 2.300 1.450 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_16


MACRO gf180mcu_osu_sc_gp9t3v3__buf_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_8 ;
  SIZE 9.050 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 2.600 1.500 2.650 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 1.100 2.250 1.500 2.300 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 5.610001 ;
    PORT
      LAYER Metal2 ;
        RECT 7.250 3.550 7.750 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 6.952500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 9.050 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 9.050 6.350 ;
        RECT 1.400 3.600 1.650 5.650 ;
        RECT 3.100 3.600 3.350 5.650 ;
        RECT 4.800 3.600 5.050 5.650 ;
        RECT 6.500 3.600 6.750 5.650 ;
        RECT 8.200 3.600 8.450 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.657500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 4.800 0.700 5.050 1.900 ;
        RECT 6.500 0.700 6.750 1.900 ;
        RECT 8.200 0.700 8.450 1.900 ;
        RECT 0.000 0.000 9.050 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.350 0.800 5.300 ;
        RECT 2.250 3.350 2.500 5.300 ;
        RECT 3.950 3.350 4.200 5.300 ;
        RECT 5.650 3.350 5.900 5.300 ;
        RECT 7.350 3.900 7.600 5.300 ;
        RECT 7.250 3.600 7.750 3.900 ;
        RECT 7.350 3.350 7.600 3.600 ;
        RECT 0.550 3.050 2.000 3.350 ;
        RECT 2.250 3.050 7.600 3.350 ;
        RECT 0.550 1.050 0.800 3.050 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 2.250 2.450 2.500 3.050 ;
        RECT 3.950 2.450 4.200 3.050 ;
        RECT 5.650 2.450 5.900 3.050 ;
        RECT 7.350 2.450 7.600 3.050 ;
        RECT 2.250 2.150 7.600 2.450 ;
        RECT 2.250 1.050 2.500 2.150 ;
        RECT 3.950 1.050 4.200 2.150 ;
        RECT 5.650 1.050 5.900 2.150 ;
        RECT 7.350 1.050 7.600 2.150 ;
      LAYER Via1 ;
        RECT 7.350 3.600 7.650 3.900 ;
        RECT 1.150 2.300 1.450 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_8


MACRO gf180mcu_osu_sc_gp9t3v3__fill_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_1 ;
  SIZE 0.900 BY 6.350 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.650 0.100 6.350 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 0.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 3.150 0.100 6.350 ;
  END
END gf180mcu_osu_sc_gp9t3v3__fill_1


MACRO gf180mcu_osu_sc_gp9t3v3__tbuf_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tbuf_1 ;
  SIZE 5.350 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.000 3.250 1.400 3.300 ;
        RECT 0.950 2.950 1.450 3.250 ;
        RECT 1.000 2.900 1.400 2.950 ;
    END
  END A
  PIN EN
    ANTENNAGATEAREA 1.020000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.750 2.250 4.250 2.650 ;
    END
  END EN
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.800 4.200 3.300 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.305000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 5.350 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 5.350 6.350 ;
        RECT 1.400 4.000 1.750 5.650 ;
        RECT 3.650 3.600 3.900 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.327500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.750 1.900 ;
        RECT 3.650 0.700 3.900 1.900 ;
        RECT 0.000 0.000 5.350 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.900 0.800 5.300 ;
        RECT 0.450 3.500 0.800 3.900 ;
        RECT 2.900 4.650 3.150 5.300 ;
        RECT 2.900 4.150 3.200 4.650 ;
        RECT 2.900 3.750 3.150 4.150 ;
        RECT 2.450 3.500 3.150 3.750 ;
        RECT 0.450 2.500 0.700 3.500 ;
        RECT 0.950 2.950 1.450 3.250 ;
        RECT 0.450 2.200 2.150 2.500 ;
        RECT 0.450 1.900 0.700 2.200 ;
        RECT 2.450 1.900 2.700 3.500 ;
        RECT 4.500 3.250 4.750 5.300 ;
        RECT 3.050 2.950 4.750 3.250 ;
        RECT 3.750 2.300 4.250 2.600 ;
        RECT 0.450 1.600 0.800 1.900 ;
        RECT 2.450 1.650 3.150 1.900 ;
        RECT 0.550 1.050 0.800 1.600 ;
        RECT 2.900 1.050 3.150 1.650 ;
        RECT 4.500 1.050 4.750 2.950 ;
      LAYER Via1 ;
        RECT 2.900 4.250 3.200 4.550 ;
        RECT 1.050 2.950 1.350 3.250 ;
        RECT 3.150 2.950 3.450 3.250 ;
        RECT 3.850 2.300 4.150 2.600 ;
      LAYER Metal2 ;
        RECT 3.050 2.900 3.550 3.300 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tbuf_1


MACRO gf180mcu_osu_sc_gp9t3v3__dlat_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dlat_1 ;
  SIZE 9.500 BY 6.350 ;
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.850 2.900 2.350 3.300 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.700 3.400 6.200 3.450 ;
        RECT 3.500 3.300 6.200 3.400 ;
        RECT 3.450 3.250 6.200 3.300 ;
        RECT 3.400 3.100 6.200 3.250 ;
        RECT 3.400 2.950 3.900 3.100 ;
        RECT 5.700 3.050 6.200 3.100 ;
        RECT 3.450 2.900 3.850 2.950 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.700 3.250 9.100 3.300 ;
        RECT 8.650 2.950 9.150 3.250 ;
        RECT 8.700 2.900 9.100 2.950 ;
    END
  END Q
  PIN VDD
    ANTENNADIFFAREA 5.167500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 9.500 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 9.500 6.350 ;
        RECT 1.450 4.400 1.700 5.650 ;
        RECT 5.350 3.850 5.600 5.650 ;
        RECT 7.800 4.300 8.050 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.020000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 0.700 1.850 1.600 ;
        RECT 5.200 0.700 5.600 1.550 ;
        RECT 7.800 0.700 8.050 1.550 ;
        RECT 0.000 0.000 9.500 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.600 2.650 0.850 5.300 ;
        RECT 3.150 4.150 3.400 5.300 ;
        RECT 1.150 3.900 3.400 4.150 ;
        RECT 6.200 4.000 6.450 5.300 ;
        RECT 1.150 3.400 1.400 3.900 ;
        RECT 6.200 3.750 6.700 4.000 ;
        RECT 1.100 3.100 1.550 3.400 ;
        RECT 0.500 2.600 0.850 2.650 ;
        RECT 0.350 2.300 0.850 2.600 ;
        RECT 0.450 2.250 0.850 2.300 ;
        RECT 0.600 1.050 0.850 2.250 ;
        RECT 1.150 2.250 1.400 3.100 ;
        RECT 1.850 2.950 2.350 3.250 ;
        RECT 2.600 3.100 3.100 3.400 ;
        RECT 2.700 2.700 3.000 3.100 ;
        RECT 3.400 2.950 3.900 3.400 ;
        RECT 5.700 3.100 6.200 3.400 ;
        RECT 4.150 2.700 4.650 2.850 ;
        RECT 2.700 2.550 4.650 2.700 ;
        RECT 2.700 2.450 4.550 2.550 ;
        RECT 5.000 2.450 5.500 2.750 ;
        RECT 2.700 2.400 4.500 2.450 ;
        RECT 1.150 2.000 2.400 2.250 ;
        RECT 2.150 1.550 2.400 2.000 ;
        RECT 4.200 2.050 4.500 2.400 ;
        RECT 6.450 2.350 6.700 3.750 ;
        RECT 6.950 3.700 7.200 5.300 ;
        RECT 6.950 3.450 8.300 3.700 ;
        RECT 7.200 2.450 7.700 2.750 ;
        RECT 6.200 2.100 6.700 2.350 ;
        RECT 8.000 2.200 8.300 3.450 ;
        RECT 6.200 2.050 6.450 2.100 ;
        RECT 4.200 1.800 6.450 2.050 ;
        RECT 3.150 1.550 3.400 1.650 ;
        RECT 2.150 1.300 3.400 1.550 ;
        RECT 3.150 1.050 3.400 1.300 ;
        RECT 6.200 1.050 6.450 1.800 ;
        RECT 6.950 1.950 8.300 2.200 ;
        RECT 8.650 3.300 8.900 5.300 ;
        RECT 8.650 3.250 9.050 3.300 ;
        RECT 8.650 2.950 9.150 3.250 ;
        RECT 8.650 2.900 9.050 2.950 ;
        RECT 6.950 1.050 7.200 1.950 ;
        RECT 8.650 1.050 8.900 2.900 ;
      LAYER Via1 ;
        RECT 0.450 2.300 0.750 2.600 ;
        RECT 1.950 2.950 2.250 3.250 ;
        RECT 3.500 2.950 3.800 3.250 ;
        RECT 5.800 3.100 6.100 3.400 ;
        RECT 5.100 2.450 5.400 2.750 ;
        RECT 7.300 2.450 7.600 2.750 ;
        RECT 8.750 2.950 9.050 3.250 ;
      LAYER Metal2 ;
        RECT 5.050 2.750 5.450 2.800 ;
        RECT 7.200 2.750 7.700 2.800 ;
        RECT 0.350 2.600 0.850 2.650 ;
        RECT 4.600 2.600 7.700 2.750 ;
        RECT 0.350 2.450 7.700 2.600 ;
        RECT 0.350 2.400 5.450 2.450 ;
        RECT 7.200 2.400 7.700 2.450 ;
        RECT 0.350 2.300 4.900 2.400 ;
        RECT 0.350 2.250 0.850 2.300 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dlat_1


MACRO gf180mcu_osu_sc_gp9t3v3__inv_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_1 ;
  SIZE 2.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.550 2.250 1.050 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 3.550 1.800 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 2.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 2.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.762500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.900 1.650 5.300 ;
        RECT 1.300 3.600 1.800 3.900 ;
        RECT 0.550 2.300 1.050 2.600 ;
        RECT 1.400 1.050 1.650 3.600 ;
      LAYER Via1 ;
        RECT 1.400 3.600 1.700 3.900 ;
        RECT 0.650 2.300 0.950 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__inv_1


MACRO gf180mcu_osu_sc_gp9t3v3__and2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__and2_1 ;
  SIZE 4.100 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.650 2.600 1.050 2.650 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 0.650 2.250 1.050 2.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.950 2.900 2.450 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.300 3.550 3.800 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.137500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 4.100 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 4.100 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.250 3.600 2.700 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.777500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.700 2.700 1.900 ;
        RECT 0.000 0.000 4.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 2.600 1.650 5.300 ;
        RECT 3.300 3.950 3.550 5.300 ;
        RECT 3.300 3.900 3.700 3.950 ;
        RECT 3.300 3.600 3.800 3.900 ;
        RECT 3.300 3.550 3.700 3.600 ;
        RECT 1.950 2.950 2.450 3.250 ;
        RECT 2.750 2.600 3.050 2.700 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 1.400 2.300 3.050 2.600 ;
        RECT 1.400 1.800 1.650 2.300 ;
        RECT 2.750 2.200 3.050 2.300 ;
        RECT 0.700 1.550 1.650 1.800 ;
        RECT 0.700 1.050 0.950 1.550 ;
        RECT 3.300 1.050 3.550 3.550 ;
      LAYER Via1 ;
        RECT 3.400 3.600 3.700 3.900 ;
        RECT 2.050 2.950 2.350 3.250 ;
        RECT 0.700 2.300 1.000 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__and2_1


MACRO gf180mcu_osu_sc_gp9t3v3__oai21_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai21_1 ;
  SIZE 4.000 BY 6.350 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 2.250 1.100 2.650 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.650 2.900 2.150 3.300 ;
    END
  END A1
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.350 2.250 2.850 2.650 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.050 3.900 3.450 3.950 ;
        RECT 3.000 3.600 3.500 3.900 ;
        RECT 3.050 3.550 3.450 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.730000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 4.000 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 4.000 6.350 ;
        RECT 0.650 3.600 0.900 5.650 ;
        RECT 3.050 4.550 3.300 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.480000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 0.700 1.600 1.500 ;
        RECT 0.000 0.000 4.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.100 3.900 2.450 5.300 ;
        RECT 2.100 3.600 3.500 3.900 ;
        RECT 3.100 3.550 3.450 3.600 ;
        RECT 1.650 2.950 2.150 3.250 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 2.350 2.300 2.850 2.600 ;
        RECT 0.500 1.750 2.550 2.000 ;
        RECT 0.500 1.050 0.750 1.750 ;
        RECT 2.200 1.050 2.550 1.750 ;
        RECT 3.150 1.050 3.400 3.550 ;
      LAYER Via1 ;
        RECT 3.100 3.600 3.400 3.900 ;
        RECT 1.750 2.950 2.050 3.250 ;
        RECT 0.700 2.300 1.000 2.600 ;
        RECT 2.450 2.300 2.750 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai21_1


MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_2 ;
  SIZE 3.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.650 2.250 1.150 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 1.600 3.900 2.000 3.950 ;
        RECT 1.550 3.600 2.050 3.900 ;
        RECT 1.600 3.550 2.000 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.460000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.300 3.600 2.550 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 0.000 0.000 3.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.900 1.650 5.300 ;
        RECT 1.400 3.600 2.050 3.900 ;
        RECT 0.650 2.300 1.150 2.600 ;
        RECT 1.400 1.050 1.650 3.600 ;
      LAYER Via1 ;
        RECT 0.750 2.300 1.050 2.600 ;
        RECT 1.650 3.600 1.950 3.900 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkinv_2


MACRO gf180mcu_osu_sc_gp9t3v3__antfill
  CLASS BLOCK ;
  ORIGIN 0 0.050 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__antfill ;
  SIZE 2.200 BY 6.350 ;
  PIN VDD
    ANTENNADIFFAREA 0.337500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.100 2.200 6.300 ;
      LAYER Metal1 ;
        RECT 0.000 5.600 2.200 6.300 ;
        RECT 1.400 3.550 1.650 5.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.337500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.050 2.200 0.650 ;
    END
  END VSS
  PIN A
    PORT
      LAYER Metal2 ;
        RECT 0.500 2.550 0.900 2.600 ;
        RECT 0.450 2.250 0.950 2.550 ;
        RECT 0.500 2.200 0.900 2.250 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.650 0.800 5.250 ;
        RECT 0.500 2.550 0.800 2.650 ;
        RECT 0.450 2.250 1.650 2.550 ;
        RECT 0.500 2.200 0.800 2.250 ;
        RECT 0.550 1.000 0.800 2.200 ;
        RECT 1.400 1.000 1.650 2.250 ;
      LAYER Via1 ;
        RECT 0.550 2.250 0.850 2.550 ;
  END
END gf180mcu_osu_sc_gp9t3v3__antfill


MACRO gf180mcu_osu_sc_gp9t3v3__xor2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__xor2_1 ;
  SIZE 6.700 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.150 2.600 1.550 2.650 ;
        RECT 1.100 2.300 1.600 2.600 ;
        RECT 1.150 2.250 1.550 2.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.150 2.600 5.550 2.650 ;
        RECT 5.100 2.300 5.600 2.600 ;
        RECT 5.150 2.250 5.550 2.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 2.167500 ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 4.600 3.450 4.650 ;
        RECT 3.100 4.200 3.500 4.600 ;
        RECT 3.150 1.850 3.450 4.200 ;
        RECT 3.050 1.450 3.550 1.850 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.557500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 6.700 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 6.700 6.350 ;
        RECT 1.400 3.900 1.650 5.650 ;
        RECT 5.000 3.900 5.250 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.622500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 5.000 0.700 5.250 1.850 ;
        RECT 0.000 0.000 6.700 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.350 0.800 5.300 ;
        RECT 3.200 4.650 3.450 5.300 ;
        RECT 3.150 4.550 3.450 4.650 ;
        RECT 3.050 4.250 3.550 4.550 ;
        RECT 2.700 3.750 4.700 4.000 ;
        RECT 2.700 3.400 3.000 3.750 ;
        RECT 4.450 3.500 4.700 3.750 ;
        RECT 5.850 3.500 6.100 5.300 ;
        RECT 0.550 3.100 2.350 3.350 ;
        RECT 2.600 3.150 3.100 3.400 ;
        RECT 0.550 1.050 0.800 3.100 ;
        RECT 2.050 2.900 2.350 3.100 ;
        RECT 3.650 2.900 3.950 3.500 ;
        RECT 4.450 3.200 6.100 3.500 ;
        RECT 4.450 2.950 4.750 3.200 ;
        RECT 2.050 2.650 3.950 2.900 ;
        RECT 4.350 2.650 4.850 2.950 ;
        RECT 1.100 2.300 1.600 2.600 ;
        RECT 5.100 2.400 5.600 2.600 ;
        RECT 2.350 2.300 5.600 2.400 ;
        RECT 2.350 2.100 5.450 2.300 ;
        RECT 3.150 1.800 3.450 1.850 ;
        RECT 3.050 1.500 3.550 1.800 ;
        RECT 3.150 1.400 3.450 1.500 ;
        RECT 3.200 1.050 3.450 1.400 ;
        RECT 5.850 1.050 6.100 3.200 ;
      LAYER Via1 ;
        RECT 3.150 4.250 3.450 4.550 ;
        RECT 1.200 2.300 1.500 2.600 ;
        RECT 5.200 2.300 5.500 2.600 ;
        RECT 3.150 1.500 3.450 1.800 ;
  END
END gf180mcu_osu_sc_gp9t3v3__xor2_1


MACRO gf180mcu_osu_sc_gp9t3v3__inv_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_2 ;
  SIZE 3.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.650 2.250 1.150 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 1.600 3.900 2.000 3.950 ;
        RECT 1.550 3.600 2.050 3.900 ;
        RECT 1.600 3.550 2.000 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.460000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.300 3.600 2.550 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 0.000 0.000 3.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.900 1.650 5.300 ;
        RECT 1.400 3.600 2.050 3.900 ;
        RECT 0.650 2.300 1.150 2.600 ;
        RECT 1.400 1.050 1.650 3.600 ;
      LAYER Via1 ;
        RECT 0.750 2.300 1.050 2.600 ;
        RECT 1.650 3.600 1.950 3.900 ;
  END
END gf180mcu_osu_sc_gp9t3v3__inv_2


MACRO gf180mcu_osu_sc_gp9t3v3__oai22_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai22_1 ;
  SIZE 5.500 BY 6.350 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.700 2.250 1.200 2.650 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.650 2.250 2.150 2.650 ;
    END
  END A1
  PIN B0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.550 2.250 3.050 2.650 ;
    END
  END B0
  PIN B1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.350 2.250 3.850 2.650 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA 1.572500 ;
    PORT
      LAYER Metal2 ;
        RECT 3.050 1.250 3.550 1.300 ;
        RECT 4.550 1.250 4.950 1.300 ;
        RECT 3.050 0.950 5.000 1.250 ;
        RECT 3.050 0.900 3.550 0.950 ;
        RECT 4.550 0.900 4.950 0.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 3.050000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 5.500 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 5.500 6.350 ;
        RECT 0.650 3.600 0.900 5.650 ;
        RECT 3.600 3.600 3.850 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.817500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 0.700 1.600 1.550 ;
        RECT 0.000 0.000 5.500 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.100 3.150 2.450 5.300 ;
        RECT 2.100 2.850 4.900 3.150 ;
        RECT 0.700 2.300 1.200 2.600 ;
        RECT 1.650 2.300 2.150 2.600 ;
        RECT 2.550 2.300 3.050 2.600 ;
        RECT 3.350 2.300 3.850 2.600 ;
        RECT 0.500 1.800 4.250 2.050 ;
        RECT 0.500 1.050 0.750 1.800 ;
        RECT 2.200 1.050 2.550 1.800 ;
        RECT 3.150 1.300 3.400 1.550 ;
        RECT 3.050 0.950 3.550 1.300 ;
        RECT 4.000 1.050 4.250 1.800 ;
        RECT 4.600 1.250 4.900 2.850 ;
        RECT 4.500 0.950 5.000 1.250 ;
      LAYER Via1 ;
        RECT 0.800 2.300 1.100 2.600 ;
        RECT 1.750 2.300 2.050 2.600 ;
        RECT 2.650 2.300 2.950 2.600 ;
        RECT 3.450 2.300 3.750 2.600 ;
        RECT 3.150 0.950 3.450 1.250 ;
        RECT 4.600 0.950 4.900 1.250 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai22_1


MACRO gf180mcu_osu_sc_gp9t3v3__dffsr_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dffsr_1 ;
  SIZE 22.100 BY 6.350 ;
  PIN D
    ANTENNAGATEAREA 0.690000 ;
    PORT
      LAYER Metal2 ;
        RECT 6.050 3.250 6.550 3.300 ;
        RECT 6.000 2.950 6.600 3.250 ;
        RECT 6.050 2.900 6.550 2.950 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.350 3.250 13.750 3.300 ;
        RECT 13.300 2.950 13.800 3.250 ;
        RECT 13.350 2.900 13.750 2.950 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.150 4.550 21.550 4.600 ;
        RECT 21.100 4.250 21.600 4.550 ;
        RECT 21.150 4.200 21.550 4.250 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 0.765000 ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 20.550 3.900 20.950 3.950 ;
        RECT 20.500 3.600 21.000 3.900 ;
        RECT 20.550 3.550 20.950 3.600 ;
    END
  END QN
  PIN S
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 18.100 3.450 18.400 3.900 ;
        RECT 18.050 3.400 18.450 3.450 ;
        RECT 18.000 3.100 18.500 3.400 ;
        RECT 18.050 3.050 18.450 3.100 ;
    END
  END S
  PIN R
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.750 3.250 1.150 3.300 ;
        RECT 0.700 2.950 1.200 3.250 ;
        RECT 0.750 2.900 1.150 2.950 ;
    END
  END R
  PIN VDD
    ANTENNADIFFAREA 12.962501 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 22.100 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 22.100 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 3.850 4.350 4.100 5.650 ;
        RECT 5.700 4.850 5.950 5.650 ;
        RECT 9.300 4.200 9.550 5.650 ;
        RECT 12.900 4.850 13.150 5.650 ;
        RECT 15.500 4.350 15.750 5.650 ;
        RECT 17.950 4.100 18.200 5.650 ;
        RECT 20.400 4.150 20.650 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 10.040001 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.300 0.700 2.550 1.500 ;
        RECT 4.550 0.700 4.800 1.550 ;
        RECT 5.700 0.700 5.950 1.600 ;
        RECT 9.300 0.700 9.550 1.500 ;
        RECT 12.900 0.700 13.150 1.800 ;
        RECT 14.800 0.700 15.050 1.900 ;
        RECT 17.050 0.700 17.300 1.500 ;
        RECT 17.950 0.700 18.200 1.900 ;
        RECT 20.400 0.700 20.650 1.700 ;
        RECT 0.000 0.000 22.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.800 2.850 1.100 3.350 ;
        RECT 1.400 2.650 1.650 5.300 ;
        RECT 1.400 2.600 1.700 2.650 ;
        RECT 1.400 2.300 1.800 2.600 ;
        RECT 1.400 2.000 1.700 2.300 ;
        RECT 2.150 2.000 2.400 5.300 ;
        RECT 3.000 4.100 3.250 5.300 ;
        RECT 4.700 4.100 4.950 5.300 ;
        RECT 7.600 4.600 8.150 5.300 ;
        RECT 3.000 3.850 4.950 4.100 ;
        RECT 5.400 4.300 8.150 4.600 ;
        RECT 5.400 3.400 5.700 4.300 ;
        RECT 10.700 3.950 11.250 5.300 ;
        RECT 12.350 4.300 12.850 4.600 ;
        RECT 12.450 4.200 12.750 4.300 ;
        RECT 13.750 4.200 14.000 5.300 ;
        RECT 13.750 3.900 14.300 4.200 ;
        RECT 6.900 3.400 13.550 3.700 ;
        RECT 3.400 3.100 3.900 3.400 ;
        RECT 4.400 3.100 5.700 3.400 ;
        RECT 5.400 2.600 5.700 3.100 ;
        RECT 6.050 2.950 6.550 3.250 ;
        RECT 6.800 3.100 7.300 3.400 ;
        RECT 2.650 2.300 3.150 2.600 ;
        RECT 5.400 2.300 6.550 2.600 ;
        RECT 10.350 2.550 10.650 3.400 ;
        RECT 13.300 3.250 13.700 3.400 ;
        RECT 11.400 2.850 11.900 3.150 ;
        RECT 13.300 2.950 13.800 3.250 ;
        RECT 3.850 2.000 5.150 2.300 ;
        RECT 1.400 1.050 1.650 2.000 ;
        RECT 2.150 1.750 4.100 2.000 ;
        RECT 3.150 1.700 4.100 1.750 ;
        RECT 6.250 1.750 6.550 2.300 ;
        RECT 7.000 2.250 7.500 2.550 ;
        RECT 9.000 2.400 9.300 2.450 ;
        RECT 8.900 2.100 9.400 2.400 ;
        RECT 10.250 2.300 10.750 2.550 ;
        RECT 11.500 2.300 11.800 2.850 ;
        RECT 12.350 2.550 12.850 2.850 ;
        RECT 14.050 2.600 14.300 3.900 ;
        RECT 14.650 4.100 14.900 5.300 ;
        RECT 16.350 4.100 16.600 5.300 ;
        RECT 14.650 3.850 16.600 4.100 ;
        RECT 17.200 4.200 17.450 5.300 ;
        RECT 18.800 4.550 19.050 5.300 ;
        RECT 18.750 4.250 19.200 4.550 ;
        RECT 17.200 3.950 17.500 4.200 ;
        RECT 14.550 2.950 15.650 3.250 ;
        RECT 15.900 2.950 16.400 3.250 ;
        RECT 13.750 2.300 14.300 2.600 ;
        RECT 11.500 2.050 14.000 2.300 ;
        RECT 14.600 2.150 15.100 2.450 ;
        RECT 3.150 1.050 3.400 1.700 ;
        RECT 6.250 1.500 8.150 1.750 ;
        RECT 7.600 1.050 8.150 1.500 ;
        RECT 10.700 1.050 11.250 1.950 ;
        RECT 13.750 1.050 14.000 2.050 ;
        RECT 15.350 2.000 15.650 2.950 ;
        RECT 17.250 2.750 17.500 3.950 ;
        RECT 18.800 3.550 19.100 4.250 ;
        RECT 19.550 3.900 19.800 5.300 ;
        RECT 21.250 4.650 21.500 5.300 ;
        RECT 21.200 4.150 21.500 4.650 ;
        RECT 19.550 3.600 21.000 3.900 ;
        RECT 20.600 3.550 20.900 3.600 ;
        RECT 18.100 3.400 18.400 3.500 ;
        RECT 18.000 3.100 18.500 3.400 ;
        RECT 18.100 3.050 18.400 3.100 ;
        RECT 19.550 2.750 20.200 2.950 ;
        RECT 17.250 2.650 20.200 2.750 ;
        RECT 16.500 2.250 17.000 2.550 ;
        RECT 17.250 2.450 19.800 2.650 ;
        RECT 17.250 2.000 17.500 2.450 ;
        RECT 20.650 2.200 20.900 3.550 ;
        RECT 15.350 1.750 17.500 2.000 ;
        RECT 18.700 1.850 19.200 2.150 ;
        RECT 19.550 1.950 20.900 2.200 ;
        RECT 16.200 1.050 16.450 1.750 ;
        RECT 18.800 1.050 19.050 1.850 ;
        RECT 19.550 1.050 19.800 1.950 ;
        RECT 21.250 1.050 21.500 4.150 ;
      LAYER Via1 ;
        RECT 0.800 2.950 1.100 3.250 ;
        RECT 10.800 4.050 11.100 4.350 ;
        RECT 12.450 4.300 12.750 4.600 ;
        RECT 3.500 3.100 3.800 3.400 ;
        RECT 4.500 3.100 4.800 3.400 ;
        RECT 6.150 2.950 6.450 3.250 ;
        RECT 2.750 2.300 3.050 2.600 ;
        RECT 13.400 2.950 13.700 3.250 ;
        RECT 4.750 2.000 5.050 2.300 ;
        RECT 7.100 2.250 7.400 2.550 ;
        RECT 9.000 2.100 9.300 2.400 ;
        RECT 11.500 2.350 11.800 2.650 ;
        RECT 12.450 2.550 12.750 2.850 ;
        RECT 18.800 4.250 19.100 4.550 ;
        RECT 14.650 2.950 14.950 3.250 ;
        RECT 16.000 2.950 16.300 3.250 ;
        RECT 14.700 2.150 15.000 2.450 ;
        RECT 10.800 1.650 11.100 1.950 ;
        RECT 21.200 4.250 21.500 4.550 ;
        RECT 20.600 3.600 20.900 3.900 ;
        RECT 18.100 3.100 18.400 3.400 ;
        RECT 16.600 2.250 16.900 2.550 ;
        RECT 19.800 2.650 20.100 2.950 ;
        RECT 18.800 1.850 19.100 2.150 ;
      LAYER Metal2 ;
        RECT 3.500 5.350 16.300 5.650 ;
        RECT 3.500 3.450 3.800 5.350 ;
        RECT 7.100 4.750 11.800 5.050 ;
        RECT 3.400 3.050 3.900 3.450 ;
        RECT 4.400 3.050 4.900 3.450 ;
        RECT 1.350 2.600 1.750 2.650 ;
        RECT 2.650 2.600 3.150 2.650 ;
        RECT 7.100 2.600 7.400 4.750 ;
        RECT 10.800 4.400 11.100 4.450 ;
        RECT 10.750 4.000 11.150 4.400 ;
        RECT 1.300 2.300 3.150 2.600 ;
        RECT 7.050 2.550 7.500 2.600 ;
        RECT 1.350 2.250 1.750 2.300 ;
        RECT 2.650 2.250 3.150 2.300 ;
        RECT 4.650 2.300 5.150 2.350 ;
        RECT 2.750 1.300 3.050 2.250 ;
        RECT 4.650 2.000 6.600 2.300 ;
        RECT 7.000 2.250 7.500 2.550 ;
        RECT 9.000 2.450 9.300 2.500 ;
        RECT 7.050 2.200 7.500 2.250 ;
        RECT 8.950 2.400 9.350 2.450 ;
        RECT 4.650 1.950 5.150 2.000 ;
        RECT 6.300 1.900 6.600 2.000 ;
        RECT 8.950 2.100 9.400 2.400 ;
        RECT 8.950 2.050 9.350 2.100 ;
        RECT 8.950 1.900 9.300 2.050 ;
        RECT 10.800 2.000 11.100 4.000 ;
        RECT 11.500 2.700 11.800 4.750 ;
        RECT 12.400 4.600 12.800 4.650 ;
        RECT 12.350 4.300 14.500 4.600 ;
        RECT 12.400 4.250 12.800 4.300 ;
        RECT 12.450 2.900 12.750 4.250 ;
        RECT 14.200 3.300 14.500 4.300 ;
        RECT 16.000 4.550 16.300 5.350 ;
        RECT 18.750 4.550 19.150 4.600 ;
        RECT 16.000 4.250 19.150 4.550 ;
        RECT 16.000 3.300 16.300 4.250 ;
        RECT 18.750 4.200 19.150 4.250 ;
        RECT 14.200 2.950 15.050 3.300 ;
        RECT 14.550 2.900 15.050 2.950 ;
        RECT 15.900 2.900 16.400 3.300 ;
        RECT 12.400 2.850 12.800 2.900 ;
        RECT 11.450 2.300 11.850 2.700 ;
        RECT 12.350 2.550 12.850 2.850 ;
        RECT 16.600 2.600 16.900 2.650 ;
        RECT 12.400 2.500 12.800 2.550 ;
        RECT 11.500 2.250 11.800 2.300 ;
        RECT 14.600 2.100 15.100 2.500 ;
        RECT 16.550 2.150 16.950 2.600 ;
        RECT 18.800 2.200 19.100 4.200 ;
        RECT 19.750 2.950 20.150 3.000 ;
        RECT 19.600 2.650 20.200 2.950 ;
        RECT 19.750 2.600 20.150 2.650 ;
        RECT 10.750 1.950 11.150 2.000 ;
        RECT 14.600 1.950 15.000 2.100 ;
        RECT 6.300 1.600 9.300 1.900 ;
        RECT 10.700 1.650 15.000 1.950 ;
        RECT 10.750 1.600 11.150 1.650 ;
        RECT 16.550 1.300 16.850 2.150 ;
        RECT 18.700 1.800 19.200 2.200 ;
        RECT 2.750 1.000 16.850 1.300 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dffsr_1


MACRO gf180mcu_osu_sc_gp9t3v3__aoi22_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__aoi22_1 ;
  SIZE 5.400 BY 6.350 ;
  PIN A0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 2.250 1.100 2.650 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.600 2.900 2.100 3.300 ;
    END
  END A1
  PIN B0
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.400 2.900 2.900 3.300 ;
    END
  END B0
  PIN B1
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.300 2.900 3.800 3.300 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 3.000 4.550 3.500 4.600 ;
        RECT 4.450 4.550 4.850 4.650 ;
        RECT 3.000 4.250 4.850 4.550 ;
        RECT 3.000 4.200 3.500 4.250 ;
        RECT 4.450 4.150 4.850 4.250 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.285000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 5.400 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 5.400 6.350 ;
        RECT 1.400 4.350 1.650 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.200000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 0.700 0.950 1.900 ;
        RECT 3.500 0.700 3.750 1.900 ;
        RECT 0.000 0.000 5.400 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.000 0.800 5.300 ;
        RECT 2.250 4.000 2.500 5.300 ;
        RECT 3.100 4.550 3.350 5.300 ;
        RECT 3.000 4.250 3.500 4.550 ;
        RECT 3.950 4.000 4.250 5.300 ;
        RECT 4.500 4.150 4.800 4.650 ;
        RECT 0.550 3.750 4.250 4.000 ;
        RECT 1.600 2.950 2.100 3.250 ;
        RECT 2.400 2.950 2.900 3.250 ;
        RECT 3.300 2.950 3.800 3.250 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 4.550 2.400 4.800 4.150 ;
        RECT 2.100 2.150 4.800 2.400 ;
        RECT 2.100 1.050 2.350 2.150 ;
      LAYER Via1 ;
        RECT 3.100 4.250 3.400 4.550 ;
        RECT 4.500 4.250 4.800 4.550 ;
        RECT 1.700 2.950 2.000 3.250 ;
        RECT 2.500 2.950 2.800 3.250 ;
        RECT 3.400 2.950 3.700 3.250 ;
        RECT 0.700 2.300 1.000 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__aoi22_1


MACRO gf180mcu_osu_sc_gp9t3v3__buf_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_1 ;
  SIZE 3.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 3.250 1.500 3.300 ;
        RECT 1.050 2.950 1.550 3.250 ;
        RECT 1.100 2.900 1.500 2.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.250 3.550 2.750 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.780000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.200 6.350 ;
        RECT 1.400 3.600 1.750 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.227500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.750 1.900 ;
        RECT 0.000 0.000 3.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.550 0.800 5.300 ;
        RECT 2.350 3.900 2.600 5.300 ;
        RECT 2.250 3.600 2.750 3.900 ;
        RECT 1.050 2.950 1.550 3.250 ;
        RECT 0.550 2.250 2.200 2.550 ;
        RECT 0.550 1.050 0.800 2.250 ;
        RECT 2.450 1.900 2.700 3.600 ;
        RECT 2.350 1.600 2.700 1.900 ;
        RECT 2.350 1.050 2.600 1.600 ;
      LAYER Via1 ;
        RECT 2.350 3.600 2.650 3.900 ;
        RECT 1.150 2.950 1.450 3.250 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_1


MACRO gf180mcu_osu_sc_gp9t3v3__nor2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__nor2_1 ;
  SIZE 3.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 2.250 1.100 2.650 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.000 2.900 2.500 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.317500 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 3.550 1.800 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.200 6.350 ;
        RECT 0.700 3.600 0.950 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 0.000 0.000 3.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.100 3.950 2.350 5.300 ;
        RECT 1.400 3.900 2.350 3.950 ;
        RECT 1.300 3.700 2.350 3.900 ;
        RECT 1.300 3.600 1.800 3.700 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 1.400 1.050 1.650 3.600 ;
        RECT 2.000 2.950 2.500 3.250 ;
      LAYER Via1 ;
        RECT 1.400 3.600 1.700 3.900 ;
        RECT 0.700 2.300 1.000 2.600 ;
        RECT 2.100 2.950 2.400 3.250 ;
  END
END gf180mcu_osu_sc_gp9t3v3__nor2_1


MACRO gf180mcu_osu_sc_gp9t3v3__fill_4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_4 ;
  SIZE 0.900 BY 6.350 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.650 0.400 6.350 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 0.400 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 3.150 0.400 6.350 ;
  END
END gf180mcu_osu_sc_gp9t3v3__fill_4


MACRO gf180mcu_osu_sc_gp9t3v3__addf_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__addf_1 ;
  SIZE 14.000 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 2.250 1.100 2.650 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.550 3.250 1.950 3.300 ;
        RECT 1.500 2.950 2.000 3.250 ;
        RECT 1.550 2.900 1.950 2.950 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA 2.295000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.600 2.600 3.000 2.650 ;
        RECT 2.550 2.300 3.050 2.600 ;
        RECT 2.600 2.250 3.000 2.300 ;
    END
  END CI
  PIN S
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.600 3.400 12.000 3.450 ;
        RECT 11.550 3.100 12.050 3.400 ;
        RECT 11.600 3.050 12.000 3.100 ;
    END
  END S
  PIN CO
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.300 3.400 13.700 3.450 ;
        RECT 13.250 3.100 13.750 3.400 ;
        RECT 13.300 3.050 13.700 3.100 ;
    END
  END CO
  PIN VDD
    ANTENNADIFFAREA 8.302501 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 14.000 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 14.000 6.350 ;
        RECT 1.400 4.800 1.650 5.650 ;
        RECT 4.800 4.800 5.050 5.650 ;
        RECT 6.500 4.800 6.750 5.650 ;
        RECT 10.750 4.800 11.000 5.650 ;
        RECT 12.350 4.800 12.600 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 6.007501 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.500 ;
        RECT 4.800 0.700 5.050 1.500 ;
        RECT 6.500 0.700 6.750 1.500 ;
        RECT 10.750 0.700 11.000 1.500 ;
        RECT 12.350 0.700 12.600 1.500 ;
        RECT 0.000 0.000 14.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 4.550 0.800 5.300 ;
        RECT 2.250 4.550 2.500 5.300 ;
        RECT 3.100 4.800 3.400 5.300 ;
        RECT 0.550 4.300 2.500 4.550 ;
        RECT 5.650 4.550 5.900 5.300 ;
        RECT 7.350 4.550 7.600 5.300 ;
        RECT 5.650 4.300 7.600 4.550 ;
        RECT 8.100 4.250 8.600 4.550 ;
        RECT 1.600 3.750 4.000 4.050 ;
        RECT 1.600 2.850 1.900 3.750 ;
        RECT 2.150 3.200 3.450 3.500 ;
        RECT 2.150 2.600 2.400 3.200 ;
        RECT 3.200 2.750 3.450 3.200 ;
        RECT 3.700 3.400 4.000 3.750 ;
        RECT 5.850 3.700 9.950 4.000 ;
        RECT 5.850 3.400 6.150 3.700 ;
        RECT 3.700 3.100 6.150 3.400 ;
        RECT 3.700 3.000 4.000 3.100 ;
        RECT 5.850 3.000 6.150 3.100 ;
        RECT 6.400 3.150 9.100 3.450 ;
        RECT 6.400 2.750 6.700 3.150 ;
        RECT 0.600 2.300 2.400 2.600 ;
        RECT 2.650 2.200 2.950 2.700 ;
        RECT 3.200 2.450 6.700 2.750 ;
        RECT 7.050 2.200 7.350 2.850 ;
        RECT 8.800 2.750 9.100 3.150 ;
        RECT 9.650 3.000 9.950 3.700 ;
        RECT 11.600 3.450 11.850 5.300 ;
        RECT 13.200 3.450 13.450 5.300 ;
        RECT 11.600 3.400 11.900 3.450 ;
        RECT 13.200 3.400 13.650 3.450 ;
        RECT 11.600 3.100 12.050 3.400 ;
        RECT 13.200 3.100 13.750 3.400 ;
        RECT 11.600 3.050 11.900 3.100 ;
        RECT 13.200 3.050 13.650 3.100 ;
        RECT 7.800 2.450 8.300 2.750 ;
        RECT 8.700 2.450 9.200 2.750 ;
        RECT 9.750 2.350 10.600 2.650 ;
        RECT 10.850 2.450 11.350 2.750 ;
        RECT 9.750 2.200 10.050 2.350 ;
        RECT 2.650 1.900 10.050 2.200 ;
        RECT 0.500 1.050 0.800 1.550 ;
        RECT 2.200 1.050 2.500 1.550 ;
        RECT 3.100 1.050 3.400 1.550 ;
        RECT 5.650 1.050 5.950 1.550 ;
        RECT 7.300 1.050 7.600 1.550 ;
        RECT 8.200 1.050 8.500 1.550 ;
        RECT 11.600 1.050 11.850 3.050 ;
        RECT 12.450 2.450 12.950 2.750 ;
        RECT 13.200 1.050 13.450 3.050 ;
      LAYER Via1 ;
        RECT 3.100 4.900 3.400 5.200 ;
        RECT 8.200 4.250 8.500 4.550 ;
        RECT 1.600 2.950 1.900 3.250 ;
        RECT 0.700 2.300 1.000 2.600 ;
        RECT 2.650 2.300 2.950 2.600 ;
        RECT 11.650 3.100 11.950 3.400 ;
        RECT 13.350 3.100 13.650 3.400 ;
        RECT 7.900 2.450 8.200 2.750 ;
        RECT 10.950 2.450 11.250 2.750 ;
        RECT 0.500 1.150 0.800 1.450 ;
        RECT 2.200 1.150 2.500 1.450 ;
        RECT 3.100 1.150 3.400 1.450 ;
        RECT 5.650 1.150 5.950 1.450 ;
        RECT 7.300 1.150 7.600 1.450 ;
        RECT 8.200 1.150 8.500 1.450 ;
        RECT 12.550 2.450 12.850 2.750 ;
      LAYER Metal2 ;
        RECT 3.100 5.250 3.400 5.300 ;
        RECT 3.050 5.200 3.450 5.250 ;
        RECT 3.000 4.900 12.850 5.200 ;
        RECT 3.050 4.850 3.450 4.900 ;
        RECT 3.750 2.750 4.050 4.900 ;
        RECT 8.150 4.550 8.550 4.600 ;
        RECT 8.100 4.250 11.250 4.550 ;
        RECT 8.150 4.200 8.550 4.250 ;
        RECT 7.850 2.750 8.250 2.800 ;
        RECT 3.750 2.450 8.300 2.750 ;
        RECT 0.500 1.500 0.800 1.550 ;
        RECT 2.200 1.500 2.500 1.550 ;
        RECT 3.100 1.500 3.400 1.550 ;
        RECT 0.450 1.450 0.850 1.500 ;
        RECT 2.150 1.450 2.550 1.500 ;
        RECT 0.450 1.150 2.550 1.450 ;
        RECT 0.450 1.100 0.850 1.150 ;
        RECT 2.150 1.100 2.550 1.150 ;
        RECT 3.050 1.450 3.450 1.500 ;
        RECT 3.750 1.450 4.050 2.450 ;
        RECT 7.850 2.400 8.250 2.450 ;
        RECT 5.650 1.500 5.950 1.550 ;
        RECT 7.300 1.500 7.600 1.550 ;
        RECT 3.050 1.150 4.050 1.450 ;
        RECT 5.600 1.450 6.000 1.500 ;
        RECT 7.250 1.450 7.650 1.500 ;
        RECT 8.150 1.450 8.550 1.500 ;
        RECT 8.850 1.450 9.150 4.250 ;
        RECT 10.950 2.800 11.250 4.250 ;
        RECT 12.550 2.800 12.850 4.900 ;
        RECT 10.900 2.400 11.300 2.800 ;
        RECT 12.500 2.750 12.900 2.800 ;
        RECT 12.450 2.450 12.950 2.750 ;
        RECT 12.500 2.400 12.900 2.450 ;
        RECT 10.950 2.350 11.250 2.400 ;
        RECT 12.550 2.350 12.850 2.400 ;
        RECT 5.600 1.150 7.650 1.450 ;
        RECT 8.100 1.150 9.150 1.450 ;
        RECT 3.050 1.100 3.450 1.150 ;
        RECT 5.600 1.100 6.000 1.150 ;
        RECT 7.250 1.100 7.650 1.150 ;
        RECT 8.150 1.100 8.550 1.150 ;
        RECT 0.500 1.050 0.800 1.100 ;
        RECT 2.200 1.050 2.500 1.100 ;
        RECT 3.100 1.050 3.400 1.100 ;
        RECT 5.650 1.050 5.950 1.100 ;
        RECT 7.300 1.050 7.600 1.100 ;
  END
END gf180mcu_osu_sc_gp9t3v3__addf_1


MACRO gf180mcu_osu_sc_gp9t3v3__ant
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__ant ;
  SIZE 2.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    ANTENNADIFFAREA 1.700000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.500 2.600 0.950 2.650 ;
        RECT 0.450 2.300 0.950 2.600 ;
        RECT 0.500 2.250 0.950 2.300 ;
    END
  END A
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 2.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 2.200 6.350 ;
        RECT 1.400 3.600 1.650 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.337500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.700 0.800 5.300 ;
        RECT 0.500 2.600 0.800 2.700 ;
        RECT 0.450 2.300 1.650 2.600 ;
        RECT 0.500 2.250 0.800 2.300 ;
        RECT 0.550 1.050 0.800 2.250 ;
        RECT 1.400 1.050 1.650 2.300 ;
      LAYER Via1 ;
        RECT 0.550 2.300 0.850 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__ant


MACRO gf180mcu_osu_sc_gp9t3v3__buf_4
  CLASS BLOCK ;
  ORIGIN 0 0.050 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_4 ;
  SIZE 5.700 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.150 2.550 1.550 2.600 ;
        RECT 1.100 2.250 1.600 2.550 ;
        RECT 1.150 2.200 1.550 2.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.805000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.900 3.500 4.400 3.900 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 4.070000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.100 5.700 6.300 ;
      LAYER Metal1 ;
        RECT 0.000 5.600 5.700 6.300 ;
        RECT 1.450 3.550 1.700 5.600 ;
        RECT 3.150 3.550 3.400 5.600 ;
        RECT 4.850 3.550 5.100 5.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.710000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 0.650 1.700 1.850 ;
        RECT 3.150 0.650 3.400 1.850 ;
        RECT 4.850 0.650 5.100 1.850 ;
        RECT 0.000 -0.050 5.700 0.650 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.600 3.300 0.850 5.250 ;
        RECT 2.300 3.300 2.550 5.250 ;
        RECT 4.000 3.850 4.250 5.250 ;
        RECT 3.900 3.550 4.400 3.850 ;
        RECT 4.000 3.300 4.250 3.550 ;
        RECT 0.600 3.000 2.050 3.300 ;
        RECT 2.300 3.000 4.250 3.300 ;
        RECT 0.600 1.000 0.850 3.000 ;
        RECT 1.100 2.250 1.600 2.550 ;
        RECT 2.300 2.400 2.550 3.000 ;
        RECT 4.000 2.400 4.250 3.000 ;
        RECT 2.300 2.100 4.250 2.400 ;
        RECT 2.300 1.000 2.550 2.100 ;
        RECT 4.000 1.000 4.250 2.100 ;
      LAYER Via1 ;
        RECT 4.000 3.550 4.300 3.850 ;
        RECT 1.200 2.250 1.500 2.550 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_4


MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_8
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_8 ;
  SIZE 8.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 6.120000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 2.250 0.900 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 5.610001 ;
    PORT
      LAYER Metal2 ;
        RECT 6.700 3.900 7.100 3.950 ;
        RECT 6.650 3.600 7.150 3.900 ;
        RECT 6.700 3.550 7.100 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 6.615000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 8.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 8.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.250 3.600 2.500 5.650 ;
        RECT 3.950 3.600 4.200 5.650 ;
        RECT 5.650 3.600 5.900 5.650 ;
        RECT 7.400 3.600 7.650 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 4.277500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 5.650 0.700 5.900 1.900 ;
        RECT 7.350 0.700 7.600 1.900 ;
        RECT 0.000 0.000 8.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.350 1.650 5.300 ;
        RECT 3.100 3.350 3.350 5.300 ;
        RECT 4.800 3.350 5.050 5.300 ;
        RECT 6.500 3.900 6.750 5.300 ;
        RECT 6.500 3.600 7.150 3.900 ;
        RECT 6.500 3.350 6.750 3.600 ;
        RECT 1.400 3.100 6.750 3.350 ;
        RECT 0.400 2.300 0.900 2.600 ;
        RECT 1.400 2.400 1.650 3.100 ;
        RECT 3.100 2.400 3.350 3.100 ;
        RECT 4.800 2.400 5.050 3.100 ;
        RECT 6.500 2.400 6.750 3.100 ;
        RECT 1.400 2.150 6.750 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
        RECT 4.800 1.050 5.050 2.150 ;
        RECT 6.500 1.050 6.750 2.150 ;
      LAYER Via1 ;
        RECT 6.750 3.600 7.050 3.900 ;
        RECT 0.500 2.300 0.800 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkinv_8


MACRO gf180mcu_osu_sc_gp9t3v3__tiel
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tiel ;
  SIZE 2.200 BY 6.350 ;
  PIN Y
    ANTENNADIFFAREA 0.425000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 1.600 1.800 2.000 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.187500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 2.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 2.200 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 0.762500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 0.000 0.000 2.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.250 1.650 5.300 ;
        RECT 1.150 3.000 1.650 3.250 ;
        RECT 1.400 1.950 1.650 2.000 ;
        RECT 1.300 1.650 1.800 1.950 ;
        RECT 1.400 1.050 1.650 1.650 ;
      LAYER Via1 ;
        RECT 1.400 1.650 1.700 1.950 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tiel


MACRO gf180mcu_osu_sc_gp9t3v3__addh_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__addh_1 ;
  SIZE 8.600 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.500 2.600 2.000 2.650 ;
        RECT 3.900 2.600 4.400 2.650 ;
        RECT 1.500 2.300 4.400 2.600 ;
        RECT 1.500 2.250 2.000 2.300 ;
        RECT 3.900 2.250 4.400 2.300 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.200 2.450 5.500 2.500 ;
        RECT 5.150 2.050 5.550 2.450 ;
        RECT 2.400 1.950 2.800 2.000 ;
        RECT 5.150 1.950 5.500 2.050 ;
        RECT 2.350 1.650 5.500 1.950 ;
        RECT 2.400 1.600 2.800 1.650 ;
    END
  END B
  PIN S
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal2 ;
        RECT 7.700 2.900 8.200 3.300 ;
    END
  END S
  PIN CO
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 3.550 0.900 3.950 ;
    END
  END CO
  PIN VDD
    ANTENNADIFFAREA 5.595000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 8.600 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 8.600 6.350 ;
        RECT 1.400 3.600 1.650 5.650 ;
        RECT 3.100 3.600 3.350 5.650 ;
        RECT 3.850 3.600 4.100 5.650 ;
        RECT 6.650 4.600 6.900 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.960000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 6.650 0.700 6.900 1.900 ;
        RECT 0.000 0.000 8.600 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.900 0.800 5.300 ;
        RECT 0.400 3.600 0.900 3.900 ;
        RECT 0.550 1.050 0.800 3.600 ;
        RECT 2.250 3.350 2.500 5.300 ;
        RECT 5.550 3.600 6.050 5.300 ;
        RECT 7.500 3.600 8.000 5.300 ;
        RECT 1.050 3.050 3.500 3.350 ;
        RECT 5.550 3.100 5.800 3.600 ;
        RECT 6.300 3.100 6.800 3.400 ;
        RECT 7.750 3.300 8.000 3.600 ;
        RECT 7.750 3.250 8.100 3.300 ;
        RECT 1.500 2.300 2.000 2.600 ;
        RECT 2.350 2.250 2.850 2.550 ;
        RECT 2.450 1.950 2.750 2.250 ;
        RECT 2.350 1.650 2.850 1.950 ;
        RECT 3.100 1.050 3.350 3.050 ;
        RECT 4.700 2.850 6.050 3.100 ;
        RECT 7.700 2.950 8.200 3.250 ;
        RECT 7.750 2.900 8.100 2.950 ;
        RECT 3.900 2.300 4.400 2.600 ;
        RECT 3.850 1.200 4.100 1.550 ;
        RECT 4.700 1.450 4.950 2.850 ;
        RECT 5.750 2.600 6.750 2.850 ;
        RECT 5.200 2.000 5.500 2.500 ;
        RECT 6.500 2.300 7.250 2.600 ;
        RECT 5.550 1.200 5.800 1.550 ;
        RECT 3.850 0.950 5.800 1.200 ;
        RECT 7.750 1.050 8.000 2.900 ;
      LAYER Via1 ;
        RECT 0.500 3.600 0.800 3.900 ;
        RECT 3.100 3.050 3.400 3.350 ;
        RECT 6.400 3.100 6.700 3.400 ;
        RECT 1.600 2.300 1.900 2.600 ;
        RECT 2.450 1.650 2.750 1.950 ;
        RECT 7.800 2.950 8.100 3.250 ;
        RECT 4.000 2.300 4.300 2.600 ;
        RECT 5.200 2.100 5.500 2.400 ;
      LAYER Metal2 ;
        RECT 3.000 3.350 3.500 3.400 ;
        RECT 6.300 3.350 6.800 3.450 ;
        RECT 3.000 3.050 6.800 3.350 ;
        RECT 3.000 3.000 3.500 3.050 ;
  END
END gf180mcu_osu_sc_gp9t3v3__addh_1


MACRO gf180mcu_osu_sc_gp9t3v3__fill_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_16 ;
  SIZE 1.600 BY 6.350 ;
  PIN VDD
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.650 1.600 6.350 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 1.600 0.700 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 0.000 3.150 1.600 6.350 ;
  END
END gf180mcu_osu_sc_gp9t3v3__fill_16


MACRO gf180mcu_osu_sc_gp9t3v3__buf_2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_2 ;
  SIZE 3.900 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 2.600 1.500 2.650 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 1.100 2.250 1.500 2.300 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal2 ;
        RECT 2.150 3.550 2.650 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.797500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.900 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.900 6.350 ;
        RECT 1.400 3.600 1.650 5.650 ;
        RECT 3.100 3.600 3.350 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.905000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.650 1.900 ;
        RECT 3.100 0.700 3.350 1.900 ;
        RECT 0.000 0.000 3.900 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.350 0.800 5.300 ;
        RECT 2.250 3.900 2.500 5.300 ;
        RECT 2.150 3.600 2.650 3.900 ;
        RECT 0.550 3.050 2.000 3.350 ;
        RECT 0.550 1.050 0.800 3.050 ;
        RECT 1.050 2.300 1.550 2.600 ;
        RECT 2.250 1.050 2.500 3.600 ;
      LAYER Via1 ;
        RECT 2.250 3.600 2.550 3.900 ;
        RECT 1.150 2.300 1.450 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_2


MACRO gf180mcu_osu_sc_gp9t3v3__dlatn_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dlatn_1 ;
  SIZE 11.300 BY 6.350 ;
  PIN D
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.850 2.900 2.350 3.300 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.750 2.900 8.250 3.300 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.500 3.250 10.900 3.300 ;
        RECT 10.450 2.950 10.950 3.250 ;
        RECT 10.500 2.900 10.900 2.950 ;
    END
  END Q
  PIN VDD
    ANTENNADIFFAREA 6.692501 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 11.300 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 11.300 6.350 ;
        RECT 1.450 4.400 1.700 5.650 ;
        RECT 5.350 3.850 5.600 5.650 ;
        RECT 8.000 3.650 8.250 5.650 ;
        RECT 9.600 4.300 9.850 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 5.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 0.700 1.850 1.600 ;
        RECT 5.200 0.700 5.600 1.550 ;
        RECT 8.000 0.700 8.250 1.900 ;
        RECT 9.600 0.700 9.850 1.550 ;
        RECT 0.000 0.000 11.300 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.600 2.650 0.850 5.300 ;
        RECT 3.150 4.150 3.400 5.300 ;
        RECT 1.150 3.900 3.400 4.150 ;
        RECT 6.200 4.000 6.450 5.300 ;
        RECT 1.150 3.400 1.400 3.900 ;
        RECT 6.200 3.750 6.700 4.000 ;
        RECT 1.100 3.100 1.550 3.400 ;
        RECT 0.500 2.600 0.850 2.650 ;
        RECT 0.350 2.300 0.850 2.600 ;
        RECT 0.450 2.250 0.850 2.300 ;
        RECT 0.600 1.050 0.850 2.250 ;
        RECT 1.150 2.250 1.400 3.100 ;
        RECT 1.850 2.950 2.350 3.250 ;
        RECT 2.600 3.100 3.100 3.400 ;
        RECT 2.700 2.700 3.000 3.100 ;
        RECT 3.400 2.950 3.900 3.400 ;
        RECT 5.700 3.100 6.200 3.400 ;
        RECT 4.150 2.700 4.650 2.850 ;
        RECT 2.700 2.550 4.650 2.700 ;
        RECT 2.700 2.450 4.550 2.550 ;
        RECT 5.000 2.450 5.500 2.750 ;
        RECT 2.700 2.400 4.500 2.450 ;
        RECT 1.150 2.000 2.400 2.250 ;
        RECT 2.150 1.550 2.400 2.000 ;
        RECT 4.200 2.050 4.500 2.400 ;
        RECT 6.450 2.350 6.700 3.750 ;
        RECT 7.150 3.400 7.400 5.300 ;
        RECT 8.750 3.700 9.000 5.300 ;
        RECT 8.750 3.450 10.100 3.700 ;
        RECT 6.950 3.100 7.450 3.400 ;
        RECT 6.200 2.100 6.700 2.350 ;
        RECT 6.200 2.050 6.450 2.100 ;
        RECT 4.200 1.800 6.450 2.050 ;
        RECT 3.150 1.550 3.400 1.650 ;
        RECT 2.150 1.300 3.400 1.550 ;
        RECT 3.150 1.050 3.400 1.300 ;
        RECT 6.200 1.050 6.450 1.800 ;
        RECT 7.150 1.050 7.400 3.100 ;
        RECT 7.750 2.950 8.250 3.250 ;
        RECT 9.000 2.450 9.500 2.750 ;
        RECT 9.800 2.200 10.100 3.450 ;
        RECT 8.750 1.950 10.100 2.200 ;
        RECT 10.450 3.300 10.700 5.300 ;
        RECT 10.450 3.250 10.850 3.300 ;
        RECT 10.450 2.950 10.950 3.250 ;
        RECT 10.450 2.900 10.850 2.950 ;
        RECT 8.750 1.050 9.000 1.950 ;
        RECT 10.450 1.050 10.700 2.900 ;
      LAYER Via1 ;
        RECT 0.450 2.300 0.750 2.600 ;
        RECT 1.950 2.950 2.250 3.250 ;
        RECT 3.500 2.950 3.800 3.250 ;
        RECT 5.800 3.100 6.100 3.400 ;
        RECT 5.100 2.450 5.400 2.750 ;
        RECT 7.050 3.100 7.350 3.400 ;
        RECT 7.850 2.950 8.150 3.250 ;
        RECT 9.100 2.450 9.400 2.750 ;
        RECT 10.550 2.950 10.850 3.250 ;
      LAYER Metal2 ;
        RECT 5.700 3.400 6.200 3.450 ;
        RECT 6.950 3.400 7.450 3.450 ;
        RECT 3.500 3.300 7.450 3.400 ;
        RECT 3.450 3.250 7.450 3.300 ;
        RECT 3.400 3.100 7.450 3.250 ;
        RECT 3.400 2.950 3.900 3.100 ;
        RECT 5.700 3.050 6.200 3.100 ;
        RECT 6.950 3.050 7.450 3.100 ;
        RECT 3.450 2.900 3.850 2.950 ;
        RECT 5.050 2.750 5.500 2.800 ;
        RECT 9.000 2.750 9.500 2.800 ;
        RECT 0.350 2.600 0.850 2.650 ;
        RECT 4.600 2.600 5.500 2.750 ;
        RECT 0.350 2.550 5.500 2.600 ;
        RECT 8.950 2.550 9.500 2.750 ;
        RECT 0.350 2.400 9.500 2.550 ;
        RECT 0.350 2.300 4.900 2.400 ;
        RECT 0.350 2.250 0.850 2.300 ;
        RECT 5.200 2.250 9.250 2.400 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dlatn_1


MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_1 ;
  SIZE 3.200 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.100 3.250 1.500 3.300 ;
        RECT 1.050 2.950 1.550 3.250 ;
        RECT 1.100 2.900 1.500 2.950 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.250 3.550 2.750 3.950 ;
        RECT 2.350 1.950 2.650 3.550 ;
        RECT 2.250 1.550 2.750 1.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 1.780000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.200 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.200 6.350 ;
        RECT 1.400 3.600 1.750 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.227500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.750 1.900 ;
        RECT 0.000 0.000 3.200 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 2.550 0.800 5.300 ;
        RECT 2.350 3.900 2.600 5.300 ;
        RECT 2.250 3.600 2.750 3.900 ;
        RECT 1.050 2.950 1.550 3.250 ;
        RECT 0.550 2.250 2.200 2.550 ;
        RECT 0.550 1.050 0.800 2.250 ;
        RECT 2.250 1.600 2.750 1.900 ;
        RECT 2.350 1.050 2.600 1.600 ;
      LAYER Via1 ;
        RECT 2.350 3.600 2.650 3.900 ;
        RECT 1.150 2.950 1.450 3.250 ;
        RECT 2.350 1.600 2.650 1.900 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_1


MACRO gf180mcu_osu_sc_gp9t3v3__tinv_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_1 ;
  SIZE 3.850 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.650 2.600 2.050 2.650 ;
        RECT 1.600 2.300 2.100 2.600 ;
        RECT 1.650 2.250 2.050 2.300 ;
    END
  END A
  PIN EN
    ANTENNAGATEAREA 1.020000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.850 2.600 1.250 2.650 ;
        RECT 0.800 2.300 1.300 2.600 ;
        RECT 0.850 2.250 1.250 2.300 ;
        RECT 0.900 1.950 1.200 2.250 ;
        RECT 2.400 2.050 2.900 2.450 ;
        RECT 2.400 1.950 2.800 2.050 ;
        RECT 0.900 1.650 2.800 1.950 ;
    END
  END EN
  PIN Y
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.800 4.200 3.300 4.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.117500 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.850 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.850 6.350 ;
        RECT 1.400 3.600 1.750 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.565000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.700 1.750 1.900 ;
        RECT 0.000 0.000 3.850 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.550 3.900 0.800 5.300 ;
        RECT 2.900 4.650 3.150 5.300 ;
        RECT 2.900 4.150 3.200 4.650 ;
        RECT 0.400 3.600 0.900 3.900 ;
        RECT 2.900 3.850 3.400 4.150 ;
        RECT 0.550 3.300 0.800 3.600 ;
        RECT 0.300 3.050 0.800 3.300 ;
        RECT 0.300 1.900 0.550 3.050 ;
        RECT 2.500 3.000 2.800 3.500 ;
        RECT 0.800 2.300 1.300 2.600 ;
        RECT 1.600 2.300 2.100 2.600 ;
        RECT 2.500 2.000 2.800 2.500 ;
        RECT 0.300 1.650 0.800 1.900 ;
        RECT 0.550 1.050 0.800 1.650 ;
        RECT 3.150 1.600 3.400 3.850 ;
        RECT 2.900 1.350 3.400 1.600 ;
        RECT 2.900 1.050 3.150 1.350 ;
      LAYER Via1 ;
        RECT 2.900 4.250 3.200 4.550 ;
        RECT 0.500 3.600 0.800 3.900 ;
        RECT 2.500 3.100 2.800 3.400 ;
        RECT 0.900 2.300 1.200 2.600 ;
        RECT 1.700 2.300 2.000 2.600 ;
        RECT 2.500 2.100 2.800 2.400 ;
      LAYER Metal2 ;
        RECT 0.400 3.900 0.900 3.950 ;
        RECT 0.400 3.600 2.000 3.900 ;
        RECT 0.400 3.550 0.900 3.600 ;
        RECT 1.700 3.400 2.000 3.600 ;
        RECT 2.400 3.400 2.900 3.450 ;
        RECT 1.700 3.100 2.900 3.400 ;
        RECT 2.400 3.050 2.900 3.100 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_1


MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_4
  CLASS BLOCK ;
  ORIGIN 0 0.050 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_4 ;
  SIZE 5.700 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.150 2.550 1.550 2.600 ;
        RECT 1.100 2.250 1.600 2.550 ;
        RECT 1.150 2.200 1.550 2.250 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.805000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.900 3.500 4.400 3.900 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 4.070000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.100 5.700 6.300 ;
      LAYER Metal1 ;
        RECT 0.000 5.600 5.700 6.300 ;
        RECT 1.450 3.550 1.700 5.600 ;
        RECT 3.150 3.550 3.400 5.600 ;
        RECT 4.850 3.550 5.100 5.600 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 2.710000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 0.650 1.700 1.850 ;
        RECT 3.150 0.650 3.400 1.850 ;
        RECT 4.850 0.650 5.100 1.850 ;
        RECT 0.000 -0.050 5.700 0.650 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.600 3.300 0.850 5.250 ;
        RECT 2.300 3.300 2.550 5.250 ;
        RECT 4.000 3.850 4.250 5.250 ;
        RECT 3.900 3.550 4.400 3.850 ;
        RECT 4.000 3.300 4.250 3.550 ;
        RECT 0.600 3.000 2.050 3.300 ;
        RECT 2.300 3.000 4.250 3.300 ;
        RECT 0.600 1.000 0.850 3.000 ;
        RECT 1.100 2.250 1.600 2.550 ;
        RECT 2.300 2.400 2.550 3.000 ;
        RECT 4.000 2.400 4.250 3.000 ;
        RECT 2.300 2.100 4.250 2.400 ;
        RECT 2.300 1.000 2.550 2.100 ;
        RECT 4.000 1.000 4.250 2.100 ;
      LAYER Via1 ;
        RECT 4.000 3.550 4.300 3.850 ;
        RECT 1.200 2.250 1.500 2.550 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_4


MACRO gf180mcu_osu_sc_gp9t3v3__nand2_1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__nand2_1 ;
  SIZE 3.100 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.600 2.250 1.100 2.650 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.000 2.900 2.500 3.300 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA 1.360000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.300 3.550 1.800 3.950 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.375000 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 3.100 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 3.100 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.250 3.600 2.500 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.100000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.700 2.350 1.900 ;
        RECT 0.000 0.000 3.100 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.900 1.650 5.300 ;
        RECT 1.300 3.600 1.800 3.900 ;
        RECT 0.600 2.300 1.100 2.600 ;
        RECT 1.400 1.850 1.650 3.600 ;
        RECT 2.000 2.950 2.500 3.250 ;
        RECT 0.700 1.600 1.650 1.850 ;
        RECT 0.700 1.050 0.950 1.600 ;
      LAYER Via1 ;
        RECT 1.400 3.600 1.700 3.900 ;
        RECT 0.700 2.300 1.000 2.600 ;
        RECT 2.100 2.950 2.400 3.250 ;
  END
END gf180mcu_osu_sc_gp9t3v3__nand2_1


MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_16 ;
  SIZE 15.000 BY 6.350 ;
  PIN A
    ANTENNAGATEAREA 12.240001 ;
    PORT
      LAYER Metal2 ;
        RECT 0.400 2.250 0.900 2.650 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 11.220001 ;
    PORT
      LAYER Metal2 ;
        RECT 13.400 3.900 13.800 3.950 ;
        RECT 13.350 3.600 13.850 3.900 ;
        RECT 13.400 3.550 13.800 3.600 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 12.380001 ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.150 15.000 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 15.000 6.350 ;
        RECT 0.550 3.600 0.800 5.650 ;
        RECT 2.250 3.600 2.500 5.650 ;
        RECT 3.950 3.600 4.200 5.650 ;
        RECT 5.650 3.600 5.900 5.650 ;
        RECT 7.350 3.600 7.600 5.650 ;
        RECT 9.050 3.600 9.300 5.650 ;
        RECT 10.750 3.600 11.000 5.650 ;
        RECT 12.450 3.600 12.700 5.650 ;
        RECT 14.150 3.600 14.400 5.650 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 8.172501 ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 2.250 0.700 2.500 1.900 ;
        RECT 3.950 0.700 4.200 1.900 ;
        RECT 5.650 0.700 5.900 1.900 ;
        RECT 7.350 0.700 7.600 1.900 ;
        RECT 9.050 0.700 9.300 1.900 ;
        RECT 10.750 0.700 11.000 1.900 ;
        RECT 12.450 0.700 12.700 1.900 ;
        RECT 14.150 0.700 14.400 1.900 ;
        RECT 0.000 0.000 15.000 0.700 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.350 1.650 5.300 ;
        RECT 3.100 3.350 3.350 5.300 ;
        RECT 4.800 3.350 5.050 5.300 ;
        RECT 6.500 3.350 6.750 5.300 ;
        RECT 8.200 3.350 8.450 5.300 ;
        RECT 9.900 3.350 10.150 5.300 ;
        RECT 11.600 3.350 11.850 5.300 ;
        RECT 13.300 3.900 13.550 5.300 ;
        RECT 13.300 3.600 13.850 3.900 ;
        RECT 13.300 3.350 13.550 3.600 ;
        RECT 1.400 3.100 13.550 3.350 ;
        RECT 0.400 2.300 0.900 2.600 ;
        RECT 1.400 2.400 1.650 3.100 ;
        RECT 3.100 2.400 3.350 3.100 ;
        RECT 4.800 2.400 5.050 3.100 ;
        RECT 6.500 2.400 6.750 3.100 ;
        RECT 8.200 2.400 8.450 3.100 ;
        RECT 9.900 2.400 10.150 3.100 ;
        RECT 11.600 2.400 11.850 3.100 ;
        RECT 13.300 2.400 13.550 3.100 ;
        RECT 1.400 2.150 13.550 2.400 ;
        RECT 1.400 1.050 1.650 2.150 ;
        RECT 3.100 1.050 3.350 2.150 ;
        RECT 4.800 1.050 5.050 2.150 ;
        RECT 6.500 1.050 6.750 2.150 ;
        RECT 8.200 1.050 8.450 2.150 ;
        RECT 9.900 1.050 10.150 2.150 ;
        RECT 11.600 1.050 11.850 2.150 ;
        RECT 13.300 1.050 13.550 2.150 ;
      LAYER Via1 ;
        RECT 13.450 3.600 13.750 3.900 ;
        RECT 0.500 2.300 0.800 2.600 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkinv_16


END LIBRARY